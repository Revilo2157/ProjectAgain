
module divider_dshift ( i_clk, i_rst, i_dividend, i_divisor, i_start, o_ready, 
        o_quotient, o_remainder, test_si1, test_so1, test_si2, test_si3, 
        test_so3, test_se );
  input [31:0] i_dividend;
  input [31:0] i_divisor;
  output [31:0] o_quotient;
  output [31:0] o_remainder;
  input i_clk, i_rst, i_start, test_si1, test_si2, test_si3, test_se;
  output o_ready, test_so1, test_so3;
  wire   ready, reg_carry, state_reg_1_0, n838, n839, n840, n843, n845, n847,
         n849, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n870, n934, n935, n936, n937, n938, n939, n944, n945,
         n946, n947, n948, n949, n977, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1113, n1124, n1125, n1126,
         n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
         n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1296, n1297, n1864,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
         n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2783, n2784, n2785, n2786, n3053, n3116,
         n3117, n3118, n3119, n3120, n3122, n3123, n3125, n3126, n3128, n3129,
         n3131, n3132, n3134, n3136, n3138, n3140, n3142, n3144, n3146, n3148,
         n3150, n3152, n3154, n3156, n3158, n3160, n3162, n3164, n3166, n3168,
         n3170, n3172, n3174, n3176, n3178, n3180, n3182, n3184, n3185, n3187,
         n3193, n3284, n3285, n4, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n60, n61, n63, n64,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n353,
         n354, n355, n356, n357, n358, n361, n364, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n443, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n636, n637, n638, n639, n640, n641,
         n642, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n756, n757, n758, n759, n760, n761, n762, n765, n769, n770,
         n771, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n841, n842, n844, n846, n848, n850, n863, n864, n865, n866, n867,
         n868, n869, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n940,
         n942, n943, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n976, n978, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1295, n1298, n1299, n1300, n1301,
         n1303, n1305, n1307, n1308, n1309, n1310, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
         n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1576, n1577, n1578, n1579, n1580, n1581, n1583, n1584, n1585, n1586,
         n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
         n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1638,
         n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
         n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
         n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
         n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
         n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
         n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1947, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1957, n1959, n1966, n1967,
         n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
         n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
         n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
         n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2957,
         n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
         n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
         n2988, n2989, n2990, n2991, n2992, n2993, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025;
  wire   [30:2] nq;
  wire   [30:0] q;
  wire   [31:0] sdata;
  wire   [5:0] state;
  wire   [31:0] reg_a;
  wire   [31:0] reg_b;
  assign test_so1 = n214;

  OAI22_X2 U1 ( .A1(n938), .A2(n581), .B1(n582), .B2(n583), .ZN(n2009) );
  XNOR2_X2 U2 ( .A(n584), .B(n585), .ZN(n582) );
  OAI22_X2 U3 ( .A1(n939), .A2(n581), .B1(n586), .B2(n583), .ZN(n2010) );
  XOR2_X2 U4 ( .A(n2335), .B(n587), .Z(n586) );
  OAI22_X2 U5 ( .A1(n935), .A2(n581), .B1(n583), .B2(n588), .ZN(n2011) );
  XOR2_X2 U6 ( .A(n589), .B(n590), .Z(n588) );
  AOI22_X2 U7 ( .A1(n591), .A2(n592), .B1(n593), .B2(n397), .ZN(n589) );
  OAI22_X2 U8 ( .A1(n937), .A2(n581), .B1(n594), .B2(n583), .ZN(n2012) );
  XOR2_X2 U9 ( .A(n595), .B(n596), .Z(n594) );
  AOI22_X2 U10 ( .A1(n585), .A2(n584), .B1(n597), .B2(n393), .ZN(n596) );
  OAI22_X2 U11 ( .A1(n936), .A2(n581), .B1(n598), .B2(n583), .ZN(n2013) );
  XNOR2_X2 U12 ( .A(n592), .B(n591), .ZN(n598) );
  NAND2_X2 U13 ( .A1(n599), .A2(n600), .ZN(n592) );
  OAI22_X2 U14 ( .A1(n934), .A2(n581), .B1(n583), .B2(n601), .ZN(n2014) );
  XOR2_X2 U15 ( .A(n602), .B(n603), .Z(n601) );
  XOR2_X2 U16 ( .A(n479), .B(n2022), .Z(n603) );
  OAI221_X2 U17 ( .B1(n599), .B2(n604), .C1(n604), .C2(n600), .A(n605), .ZN(
        n602) );
  AOI22_X2 U18 ( .A1(n606), .A2(n590), .B1(n2335), .B2(n454), .ZN(n605) );
  OAI22_X2 U21 ( .A1(n2022), .A2(n587), .B1(n939), .B2(n607), .ZN(n584) );
  XOR2_X2 U22 ( .A(n394), .B(n607), .Z(n587) );
  XNOR2_X2 U23 ( .A(n3116), .B(n2022), .ZN(n607) );
  XNOR2_X2 U24 ( .A(n938), .B(n597), .ZN(n585) );
  NAND2_X2 U25 ( .A1(n591), .A2(n590), .ZN(n604) );
  XOR2_X2 U26 ( .A(n935), .B(n2022), .Z(n590) );
  XOR2_X2 U27 ( .A(n936), .B(n236), .Z(n591) );
  XOR2_X2 U28 ( .A(n3119), .B(n2022), .Z(n593) );
  AOI22_X2 U29 ( .A1(n396), .A2(n608), .B1(n595), .B2(n609), .ZN(n599) );
  AND2_X2 U30 ( .A1(n597), .A2(n393), .ZN(n609) );
  XNOR2_X2 U31 ( .A(n3117), .B(n2335), .ZN(n597) );
  XNOR2_X2 U32 ( .A(n937), .B(n608), .ZN(n595) );
  XOR2_X2 U33 ( .A(n3118), .B(n2022), .Z(n608) );
  OAI211_X2 U35 ( .C1(n611), .C2(n612), .A(n613), .B(n68), .ZN(n581) );
  AOI22_X2 U36 ( .A1(n2434), .A2(n3123), .B1(n615), .B2(n2431), .ZN(n614) );
  AOI22_X2 U37 ( .A1(n2434), .A2(n3126), .B1(n618), .B2(n2431), .ZN(n617) );
  AOI22_X2 U38 ( .A1(n2434), .A2(n3129), .B1(n620), .B2(n2431), .ZN(n619) );
  AOI22_X2 U39 ( .A1(n2434), .A2(n3132), .B1(n2432), .B2(n622), .ZN(n621) );
  OAI22_X2 U40 ( .A1(n3185), .A2(n2432), .B1(n2334), .B2(n2434), .ZN(n2015) );
  AOI22_X2 U41 ( .A1(n2434), .A2(n3053), .B1(n2432), .B2(n624), .ZN(n623) );
  AOI22_X2 U42 ( .A1(n2434), .A2(n3120), .B1(n626), .B2(n2431), .ZN(n625) );
  OAI22_X2 U45 ( .A1(n2434), .A2(n322), .B1(n2004), .B2(n634), .ZN(n632) );
  AOI22_X2 U47 ( .A1(n641), .A2(n642), .B1(n2338), .B2(n644), .ZN(n628) );
  OAI22_X2 U50 ( .A1(n2434), .A2(n339), .B1(n2001), .B2(n2337), .ZN(n648) );
  AOI22_X2 U52 ( .A1(n641), .A2(n652), .B1(n2338), .B2(n653), .ZN(n645) );
  OAI22_X2 U55 ( .A1(n2435), .A2(n338), .B1(n2005), .B2(n2336), .ZN(n657) );
  AOI22_X2 U57 ( .A1(n641), .A2(n660), .B1(n2338), .B2(n661), .ZN(n654) );
  OAI22_X2 U61 ( .A1(n2434), .A2(n337), .B1(n2006), .B2(n634), .ZN(n665) );
  AOI22_X2 U64 ( .A1(n641), .A2(n673), .B1(n2338), .B2(n674), .ZN(n662) );
  NAND2_X2 U65 ( .A1(n675), .A2(n676), .ZN(n995) );
  AOI221_X2 U66 ( .B1(n2339), .B2(n640), .C1(n641), .C2(n636), .A(n677), .ZN(
        n676) );
  AOI221_X2 U68 ( .B1(sdata[15]), .B2(n2430), .C1(i_dividend[15]), .C2(n2426), 
        .A(n679), .ZN(n675) );
  OAI22_X2 U69 ( .A1(n2002), .A2(n2337), .B1(n435), .B2(n2024), .ZN(n679) );
  OAI221_X2 U70 ( .B1(n2434), .B2(n335), .C1(n2428), .C2(n548), .A(n680), .ZN(
        n994) );
  AOI221_X2 U71 ( .B1(n42), .B2(n447), .C1(n681), .C2(n682), .A(n61), .ZN(n680) );
  NAND2_X2 U72 ( .A1(n683), .A2(n684), .ZN(n993) );
  AOI221_X2 U73 ( .B1(n2339), .B2(n659), .C1(n641), .C2(n658), .A(n685), .ZN(
        n684) );
  AOI221_X2 U75 ( .B1(sdata[17]), .B2(n2430), .C1(i_dividend[17]), .C2(n2426), 
        .A(n687), .ZN(n683) );
  OAI22_X2 U76 ( .A1(n2003), .A2(n2336), .B1(n423), .B2(n2024), .ZN(n687) );
  OAI211_X2 U77 ( .C1(n2429), .C2(n547), .A(n688), .B(n689), .ZN(n992) );
  AOI221_X2 U78 ( .B1(n2339), .B2(n671), .C1(n681), .C2(n690), .A(n691), .ZN(
        n689) );
  AOI22_X2 U80 ( .A1(n42), .A2(n446), .B1(sdata[18]), .B2(n2431), .ZN(n688) );
  NAND2_X2 U81 ( .A1(n692), .A2(n693), .ZN(n991) );
  AOI221_X2 U82 ( .B1(n694), .B2(n681), .C1(n641), .C2(n640), .A(n695), .ZN(
        n693) );
  AOI221_X2 U84 ( .B1(sdata[19]), .B2(n2430), .C1(i_dividend[19]), .C2(n2426), 
        .A(n696), .ZN(n692) );
  OAI22_X2 U85 ( .A1(n1982), .A2(n634), .B1(n432), .B2(n2024), .ZN(n696) );
  OAI221_X2 U86 ( .B1(n2434), .B2(n378), .C1(n2428), .C2(n546), .A(n697), .ZN(
        n990) );
  AOI221_X2 U87 ( .B1(n42), .B2(n474), .C1(n681), .C2(n698), .A(n61), .ZN(n697) );
  OAI221_X2 U88 ( .B1(n2434), .B2(n377), .C1(n2428), .C2(n545), .A(n699), .ZN(
        n989) );
  AOI221_X2 U89 ( .B1(n42), .B2(n465), .C1(n681), .C2(n700), .A(n61), .ZN(n699) );
  OAI221_X2 U90 ( .B1(n2434), .B2(n376), .C1(n2428), .C2(n544), .A(n701), .ZN(
        n988) );
  AOI221_X2 U91 ( .B1(n42), .B2(n464), .C1(n681), .C2(n702), .A(n61), .ZN(n701) );
  OAI211_X2 U92 ( .C1(n1993), .C2(n2336), .A(n703), .B(n704), .ZN(n987) );
  AOI221_X2 U93 ( .B1(sdata[23]), .B2(n2430), .C1(i_dividend[23]), .C2(n2426), 
        .A(n60), .ZN(n704) );
  AOI22_X2 U94 ( .A1(n641), .A2(n638), .B1(n2338), .B2(n640), .ZN(n703) );
  OAI211_X2 U95 ( .C1(n1994), .C2(n634), .A(n705), .B(n706), .ZN(n986) );
  AOI221_X2 U96 ( .B1(sdata[24]), .B2(n2430), .C1(i_dividend[24]), .C2(n2426), 
        .A(n60), .ZN(n706) );
  AOI22_X2 U97 ( .A1(n641), .A2(n650), .B1(n2338), .B2(n651), .ZN(n705) );
  OAI211_X2 U98 ( .C1(n1995), .C2(n2337), .A(n707), .B(n708), .ZN(n985) );
  AOI221_X2 U99 ( .B1(sdata[25]), .B2(n2430), .C1(i_dividend[25]), .C2(n2426), 
        .A(n60), .ZN(n708) );
  AOI22_X2 U100 ( .A1(n641), .A2(n440), .B1(n2338), .B2(n659), .ZN(n707) );
  OAI211_X2 U101 ( .C1(n1996), .C2(n2336), .A(n709), .B(n710), .ZN(n984) );
  AOI221_X2 U102 ( .B1(n2430), .B2(sdata[26]), .C1(i_dividend[26]), .C2(n2426), 
        .A(n60), .ZN(n710) );
  AOI22_X2 U104 ( .A1(n641), .A2(n670), .B1(n2338), .B2(n671), .ZN(n709) );
  OAI211_X2 U105 ( .C1(n2429), .C2(n543), .A(n713), .B(n714), .ZN(n983) );
  OAI211_X2 U107 ( .C1(n2429), .C2(n542), .A(n713), .B(n715), .ZN(n982) );
  OAI211_X2 U109 ( .C1(n2429), .C2(n541), .A(n713), .B(n716), .ZN(n981) );
  OAI211_X2 U111 ( .C1(n2429), .C2(n540), .A(n713), .B(n717), .ZN(n980) );
  NAND2_X2 U116 ( .A1(n672), .A2(n455), .ZN(n667) );
  OAI221_X2 U117 ( .B1(n2334), .B2(n2434), .C1(n2428), .C2(n539), .A(n720), 
        .ZN(n979) );
  OAI22_X2 U120 ( .A1(n2431), .A2(n165), .B1(n2435), .B2(n723), .ZN(n862) );
  OAI22_X2 U121 ( .A1(n2431), .A2(n164), .B1(n2435), .B2(n724), .ZN(n861) );
  OAI22_X2 U122 ( .A1(n2431), .A2(n166), .B1(n2435), .B2(n725), .ZN(n860) );
  OAI22_X2 U123 ( .A1(n2431), .A2(n167), .B1(n2435), .B2(n726), .ZN(n859) );
  OAI22_X2 U124 ( .A1(n2431), .A2(n150), .B1(n2435), .B2(n727), .ZN(n858) );
  OAI22_X2 U125 ( .A1(n2431), .A2(n147), .B1(n2435), .B2(n728), .ZN(n857) );
  OAI22_X2 U126 ( .A1(n2431), .A2(n146), .B1(n2435), .B2(n729), .ZN(n856) );
  OAI22_X2 U127 ( .A1(n2431), .A2(n145), .B1(n2435), .B2(n730), .ZN(n855) );
  OAI22_X2 U128 ( .A1(n2431), .A2(n149), .B1(n2435), .B2(n731), .ZN(n854) );
  OAI22_X2 U129 ( .A1(n2432), .A2(n144), .B1(n2435), .B2(n732), .ZN(n853) );
  OAI22_X2 U130 ( .A1(n2432), .A2(n148), .B1(n2435), .B2(n733), .ZN(n852) );
  OAI22_X2 U131 ( .A1(n2432), .A2(n162), .B1(n2435), .B2(n734), .ZN(n851) );
  AOI22_X2 U132 ( .A1(n2434), .A2(n1949), .B1(n2432), .B2(n736), .ZN(n735) );
  OAI22_X2 U133 ( .A1(n2432), .A2(n161), .B1(n2435), .B2(n299), .ZN(n849) );
  AOI22_X2 U134 ( .A1(n2434), .A2(n1947), .B1(n2432), .B2(n739), .ZN(n738) );
  OAI22_X2 U135 ( .A1(n2432), .A2(n159), .B1(n2435), .B2(n314), .ZN(n847) );
  AOI22_X2 U136 ( .A1(n2434), .A2(n1959), .B1(n2432), .B2(n742), .ZN(n741) );
  OAI22_X2 U137 ( .A1(n2432), .A2(n152), .B1(n2435), .B2(n317), .ZN(n845) );
  AOI22_X2 U138 ( .A1(n2434), .A2(n1957), .B1(n2432), .B2(n745), .ZN(n744) );
  OAI22_X2 U139 ( .A1(n2432), .A2(n157), .B1(n2435), .B2(n323), .ZN(n843) );
  AOI22_X2 U140 ( .A1(n2434), .A2(n1967), .B1(n2432), .B2(n748), .ZN(n747) );
  AOI22_X2 U141 ( .A1(n2434), .A2(n1966), .B1(n2432), .B2(n750), .ZN(n749) );
  OAI22_X2 U142 ( .A1(n2432), .A2(n168), .B1(n2435), .B2(n751), .ZN(n840) );
  OAI22_X2 U143 ( .A1(n2432), .A2(n155), .B1(n2435), .B2(n752), .ZN(n839) );
  OAI22_X2 U144 ( .A1(n2432), .A2(n154), .B1(n2435), .B2(n753), .ZN(n838) );
  OAI22_X2 U145 ( .A1(n3119), .A2(n754), .B1(n101), .B2(n172), .ZN(n2786) );
  OAI22_X2 U146 ( .A1(n3118), .A2(n754), .B1(n101), .B2(n173), .ZN(n2785) );
  OAI22_X2 U147 ( .A1(n3117), .A2(n754), .B1(n101), .B2(n174), .ZN(n2784) );
  OAI22_X2 U148 ( .A1(n3116), .A2(n754), .B1(n101), .B2(n175), .ZN(n2783) );
  OAI22_X2 U149 ( .A1(n2419), .A2(n169), .B1(n2435), .B2(n756), .ZN(n1864) );
  OAI221_X2 U150 ( .B1(n2414), .B2(n154), .C1(n2418), .C2(n538), .A(n758), 
        .ZN(n1297) );
  AOI221_X2 U151 ( .B1(n2420), .B2(n456), .C1(q[30]), .C2(n759), .A(n760), 
        .ZN(n758) );
  NOR4_X2 U152 ( .A1(q[30]), .A2(n2442), .A3(n761), .A4(n176), .ZN(n760) );
  OAI221_X2 U154 ( .B1(n2412), .B2(n549), .C1(n2334), .C2(n2407), .A(n765), 
        .ZN(n1296) );
  OAI211_X2 U156 ( .C1(n110), .C2(n2418), .A(n754), .B(n2429), .ZN(n1293) );
  OAI211_X2 U157 ( .C1(n2419), .C2(n281), .A(n770), .B(n771), .ZN(n1292) );
  AOI22_X2 U159 ( .A1(n2421), .A2(n466), .B1(n2413), .B2(n3053), .ZN(n770) );
  NAND2_X2 U160 ( .A1(n774), .A2(n775), .ZN(n1291) );
  AOI221_X2 U161 ( .B1(n40), .B2(n441), .C1(q[1]), .C2(n36), .A(n776), .ZN(
        n775) );
  NAND2_X2 U164 ( .A1(n778), .A2(n779), .ZN(n1290) );
  AOI221_X2 U165 ( .B1(n40), .B2(n414), .C1(q[2]), .C2(n780), .A(n781), .ZN(
        n779) );
  NOR4_X2 U166 ( .A1(q[2]), .A2(n398), .A3(n195), .A4(n2442), .ZN(n781) );
  NAND2_X2 U170 ( .A1(n782), .A2(n35), .ZN(n1289) );
  OAI221_X2 U171 ( .B1(n756), .B2(n946), .C1(n193), .C2(n784), .A(n785), .ZN(
        n783) );
  OR3_X2 U172 ( .A1(n2442), .A2(q[3]), .A3(n786), .ZN(n785) );
  NAND2_X2 U174 ( .A1(n787), .A2(n788), .ZN(n1288) );
  AOI221_X2 U175 ( .B1(n40), .B2(n406), .C1(q[4]), .C2(n789), .A(n790), .ZN(
        n788) );
  NOR4_X2 U176 ( .A1(q[4]), .A2(n786), .A3(n193), .A4(n2442), .ZN(n790) );
  NAND2_X2 U180 ( .A1(n791), .A2(n792), .ZN(n1287) );
  AOI221_X2 U181 ( .B1(n40), .B2(n401), .C1(q[5]), .C2(n34), .A(n793), .ZN(
        n792) );
  OAI221_X2 U184 ( .B1(n2414), .B2(n165), .C1(n2418), .C2(n487), .A(n796), 
        .ZN(n1286) );
  AOI221_X2 U185 ( .B1(n2420), .B2(n470), .C1(q[6]), .C2(n797), .A(n798), .ZN(
        n796) );
  NOR4_X2 U186 ( .A1(q[6]), .A2(n794), .A3(n196), .A4(n2442), .ZN(n798) );
  OAI221_X2 U189 ( .B1(n2414), .B2(n164), .C1(n2418), .C2(n486), .A(n799), 
        .ZN(n1285) );
  AOI221_X2 U190 ( .B1(n2420), .B2(n469), .C1(q[7]), .C2(n33), .A(n800), .ZN(
        n799) );
  OAI221_X2 U192 ( .B1(n2414), .B2(n166), .C1(n2418), .C2(n484), .A(n803), 
        .ZN(n1284) );
  AOI221_X2 U193 ( .B1(n2420), .B2(n468), .C1(q[8]), .C2(n804), .A(n805), .ZN(
        n803) );
  NOR4_X2 U194 ( .A1(q[8]), .A2(n801), .A3(n190), .A4(n2442), .ZN(n805) );
  OAI221_X2 U197 ( .B1(n2414), .B2(n167), .C1(n2418), .C2(n483), .A(n806), 
        .ZN(n1283) );
  AOI221_X2 U198 ( .B1(n2420), .B2(n467), .C1(q[9]), .C2(n32), .A(n807), .ZN(
        n806) );
  OAI221_X2 U200 ( .B1(n2414), .B2(n150), .C1(n2419), .C2(n488), .A(n810), 
        .ZN(n1282) );
  AOI221_X2 U201 ( .B1(n2420), .B2(n476), .C1(q[10]), .C2(n811), .A(n812), 
        .ZN(n810) );
  NOR4_X2 U202 ( .A1(q[10]), .A2(n808), .A3(n199), .A4(n2442), .ZN(n812) );
  OAI221_X2 U205 ( .B1(n2414), .B2(n147), .C1(n2418), .C2(n480), .A(n813), 
        .ZN(n1281) );
  AOI221_X2 U206 ( .B1(n2420), .B2(n450), .C1(q[11]), .C2(n31), .A(n814), .ZN(
        n813) );
  OAI221_X2 U208 ( .B1(n2414), .B2(n146), .C1(n2418), .C2(n489), .A(n817), 
        .ZN(n1280) );
  AOI221_X2 U209 ( .B1(n2420), .B2(n453), .C1(q[12]), .C2(n818), .A(n819), 
        .ZN(n817) );
  NOR4_X2 U210 ( .A1(q[12]), .A2(n815), .A3(n197), .A4(n2442), .ZN(n819) );
  OAI221_X2 U213 ( .B1(n2414), .B2(n145), .C1(n2418), .C2(n493), .A(n820), 
        .ZN(n1279) );
  AOI221_X2 U214 ( .B1(n2420), .B2(n449), .C1(q[13]), .C2(n30), .A(n821), .ZN(
        n820) );
  OAI221_X2 U216 ( .B1(n2414), .B2(n149), .C1(n2418), .C2(n499), .A(n824), 
        .ZN(n1278) );
  AOI221_X2 U217 ( .B1(n2421), .B2(n448), .C1(q[14]), .C2(n825), .A(n826), 
        .ZN(n824) );
  NOR4_X2 U218 ( .A1(q[14]), .A2(n822), .A3(n211), .A4(n2442), .ZN(n826) );
  OAI221_X2 U221 ( .B1(n2414), .B2(n144), .C1(n2418), .C2(n502), .A(n827), 
        .ZN(n1277) );
  AOI221_X2 U222 ( .B1(n2421), .B2(n452), .C1(q[15]), .C2(n29), .A(n828), .ZN(
        n827) );
  OAI221_X2 U224 ( .B1(n2414), .B2(n148), .C1(n2418), .C2(n505), .A(n831), 
        .ZN(n1276) );
  AOI221_X2 U225 ( .B1(n2421), .B2(n447), .C1(q[16]), .C2(n832), .A(n833), 
        .ZN(n831) );
  NOR4_X2 U226 ( .A1(q[16]), .A2(n829), .A3(n209), .A4(n2442), .ZN(n833) );
  OAI221_X2 U229 ( .B1(n2414), .B2(n162), .C1(n2419), .C2(n510), .A(n834), 
        .ZN(n1275) );
  AOI221_X2 U230 ( .B1(n2421), .B2(n451), .C1(q[17]), .C2(n28), .A(n835), .ZN(
        n834) );
  OAI221_X2 U232 ( .B1(n2414), .B2(n163), .C1(n2419), .C2(n513), .A(n841), 
        .ZN(n1274) );
  AOI221_X2 U233 ( .B1(n2421), .B2(n446), .C1(q[18]), .C2(n842), .A(n844), 
        .ZN(n841) );
  NOR4_X2 U234 ( .A1(q[18]), .A2(n836), .A3(n207), .A4(n2442), .ZN(n844) );
  OAI221_X2 U237 ( .B1(n757), .B2(n161), .C1(n2419), .C2(n511), .A(n846), .ZN(
        n1273) );
  AOI221_X2 U238 ( .B1(n2421), .B2(n475), .C1(q[19]), .C2(n27), .A(n848), .ZN(
        n846) );
  OAI221_X2 U240 ( .B1(n757), .B2(n160), .C1(n2419), .C2(n514), .A(n864), .ZN(
        n1272) );
  AOI221_X2 U241 ( .B1(n2421), .B2(n474), .C1(q[20]), .C2(n865), .A(n866), 
        .ZN(n864) );
  NOR4_X2 U242 ( .A1(q[20]), .A2(n850), .A3(n205), .A4(n2442), .ZN(n866) );
  OAI221_X2 U245 ( .B1(n2414), .B2(n159), .C1(n2419), .C2(n517), .A(n867), 
        .ZN(n1271) );
  AOI221_X2 U246 ( .B1(n2421), .B2(n465), .C1(q[21]), .C2(n26), .A(n868), .ZN(
        n867) );
  OAI221_X2 U248 ( .B1(n757), .B2(n153), .C1(n2419), .C2(n518), .A(n872), .ZN(
        n1270) );
  AOI221_X2 U249 ( .B1(n2421), .B2(n464), .C1(q[22]), .C2(n873), .A(n874), 
        .ZN(n872) );
  NOR4_X2 U250 ( .A1(q[22]), .A2(n869), .A3(n203), .A4(n2442), .ZN(n874) );
  OAI221_X2 U253 ( .B1(n757), .B2(n152), .C1(n2419), .C2(n519), .A(n875), .ZN(
        n1269) );
  AOI221_X2 U254 ( .B1(n2421), .B2(n463), .C1(q[23]), .C2(n25), .A(n876), .ZN(
        n875) );
  OAI221_X2 U256 ( .B1(n757), .B2(n158), .C1(n2419), .C2(n522), .A(n879), .ZN(
        n1268) );
  AOI221_X2 U257 ( .B1(n2421), .B2(n462), .C1(q[24]), .C2(n880), .A(n881), 
        .ZN(n879) );
  NOR4_X2 U258 ( .A1(q[24]), .A2(n877), .A3(n201), .A4(n2442), .ZN(n881) );
  OAI221_X2 U261 ( .B1(n2414), .B2(n157), .C1(n2419), .C2(n524), .A(n882), 
        .ZN(n1267) );
  AOI221_X2 U262 ( .B1(n2421), .B2(n461), .C1(q[25]), .C2(n24), .A(n883), .ZN(
        n882) );
  OAI221_X2 U264 ( .B1(n757), .B2(n151), .C1(n2419), .C2(n525), .A(n886), .ZN(
        n1266) );
  AOI221_X2 U265 ( .B1(n2421), .B2(n460), .C1(q[26]), .C2(n887), .A(n888), 
        .ZN(n886) );
  NOR4_X2 U266 ( .A1(q[26]), .A2(n884), .A3(n180), .A4(n2442), .ZN(n888) );
  OAI221_X2 U269 ( .B1(n757), .B2(n156), .C1(n2419), .C2(n529), .A(n889), .ZN(
        n1265) );
  AOI221_X2 U270 ( .B1(n2421), .B2(n459), .C1(q[27]), .C2(n23), .A(n890), .ZN(
        n889) );
  OAI221_X2 U272 ( .B1(n2414), .B2(n168), .C1(n2419), .C2(n531), .A(n893), 
        .ZN(n1264) );
  AOI221_X2 U273 ( .B1(n2420), .B2(n458), .C1(q[28]), .C2(n894), .A(n895), 
        .ZN(n893) );
  NOR4_X2 U274 ( .A1(q[28]), .A2(n891), .A3(n178), .A4(n2442), .ZN(n895) );
  OAI221_X2 U277 ( .B1(n2414), .B2(n155), .C1(n2419), .C2(n537), .A(n896), 
        .ZN(n1263) );
  AOI221_X2 U278 ( .B1(n2421), .B2(n457), .C1(q[29]), .C2(n22), .A(n897), .ZN(
        n896) );
  OR3_X2 U283 ( .A1(n178), .A2(n891), .A3(n177), .ZN(n761) );
  OR3_X2 U284 ( .A1(n180), .A2(n884), .A3(n179), .ZN(n891) );
  OR3_X2 U285 ( .A1(n201), .A2(n877), .A3(n181), .ZN(n884) );
  OR3_X2 U286 ( .A1(n203), .A2(n869), .A3(n202), .ZN(n877) );
  OR3_X2 U287 ( .A1(n205), .A2(n850), .A3(n204), .ZN(n869) );
  OR3_X2 U288 ( .A1(n207), .A2(n836), .A3(n206), .ZN(n850) );
  OR3_X2 U289 ( .A1(n209), .A2(n829), .A3(n208), .ZN(n836) );
  OR3_X2 U290 ( .A1(n211), .A2(n822), .A3(n210), .ZN(n829) );
  OR3_X2 U291 ( .A1(n197), .A2(n815), .A3(n212), .ZN(n822) );
  OR3_X2 U292 ( .A1(n198), .A2(n808), .A3(n199), .ZN(n815) );
  OR3_X2 U293 ( .A1(n190), .A2(n801), .A3(n200), .ZN(n808) );
  OR3_X2 U294 ( .A1(n196), .A2(n794), .A3(n191), .ZN(n801) );
  OR3_X2 U295 ( .A1(n193), .A2(n786), .A3(n192), .ZN(n794) );
  OAI22_X2 U297 ( .A1(n2396), .A2(n2637), .B1(n900), .B2(n901), .ZN(n1262) );
  OAI22_X2 U298 ( .A1(n2396), .A2(n2638), .B1(n901), .B2(n280), .ZN(n1261) );
  OAI22_X2 U299 ( .A1(n2396), .A2(n2639), .B1(n901), .B2(n278), .ZN(n1260) );
  OAI22_X2 U300 ( .A1(n2396), .A2(n2640), .B1(n901), .B2(n902), .ZN(n1259) );
  OAI22_X2 U301 ( .A1(n2396), .A2(n2641), .B1(n901), .B2(n903), .ZN(n1258) );
  OAI22_X2 U302 ( .A1(n2396), .A2(n2642), .B1(n901), .B2(n271), .ZN(n1257) );
  OAI22_X2 U303 ( .A1(n2396), .A2(n2643), .B1(n901), .B2(n270), .ZN(n1256) );
  OAI22_X2 U304 ( .A1(n2396), .A2(n2644), .B1(n901), .B2(n904), .ZN(n1255) );
  OAI22_X2 U305 ( .A1(n2396), .A2(n2645), .B1(n2395), .B2(n905), .ZN(n1254) );
  OAI22_X2 U306 ( .A1(n2396), .A2(n2646), .B1(n901), .B2(n906), .ZN(n1253) );
  OAI22_X2 U307 ( .A1(n2396), .A2(n2647), .B1(n901), .B2(n907), .ZN(n1252) );
  OAI22_X2 U308 ( .A1(n2396), .A2(n2648), .B1(n901), .B2(n259), .ZN(n1251) );
  OAI22_X2 U309 ( .A1(n2396), .A2(n2649), .B1(n901), .B2(n908), .ZN(n1250) );
  OAI22_X2 U310 ( .A1(n2396), .A2(n2650), .B1(n2395), .B2(n245), .ZN(n1249) );
  OAI22_X2 U311 ( .A1(n2396), .A2(n2651), .B1(n2395), .B2(n244), .ZN(n1248) );
  OAI22_X2 U312 ( .A1(n2396), .A2(n2652), .B1(n2395), .B2(n266), .ZN(n1247) );
  OAI22_X2 U313 ( .A1(n2396), .A2(n2653), .B1(n2395), .B2(n265), .ZN(n1246) );
  OAI22_X2 U314 ( .A1(n2396), .A2(n2654), .B1(n2395), .B2(n909), .ZN(n1245) );
  OAI22_X2 U315 ( .A1(n2396), .A2(n2655), .B1(n2395), .B2(n254), .ZN(n1244) );
  OAI22_X2 U316 ( .A1(n2396), .A2(n2656), .B1(n2395), .B2(n910), .ZN(n1243) );
  OAI22_X2 U317 ( .A1(n2396), .A2(n2657), .B1(n2395), .B2(n911), .ZN(n1242) );
  OAI22_X2 U318 ( .A1(n2396), .A2(n2658), .B1(n2395), .B2(n247), .ZN(n1241) );
  OAI22_X2 U319 ( .A1(n2397), .A2(n2659), .B1(n2395), .B2(n246), .ZN(n1240) );
  OAI22_X2 U320 ( .A1(n2397), .A2(n2660), .B1(n2395), .B2(n264), .ZN(n1239) );
  OAI22_X2 U321 ( .A1(n2397), .A2(n2661), .B1(n2395), .B2(n263), .ZN(n1238) );
  OAI22_X2 U322 ( .A1(n2397), .A2(n2662), .B1(n2395), .B2(n912), .ZN(n1237) );
  OAI22_X2 U323 ( .A1(n2397), .A2(n2663), .B1(n2395), .B2(n249), .ZN(n1236) );
  OAI22_X2 U324 ( .A1(n2397), .A2(n2664), .B1(n2395), .B2(n257), .ZN(n1235) );
  OAI22_X2 U325 ( .A1(n2397), .A2(n2665), .B1(n2395), .B2(n256), .ZN(n1234) );
  OAI22_X2 U326 ( .A1(n2397), .A2(n2666), .B1(n2395), .B2(n243), .ZN(n1233) );
  OAI22_X2 U327 ( .A1(n2397), .A2(n2667), .B1(n2395), .B2(n242), .ZN(n1232) );
  OAI22_X2 U328 ( .A1(n2396), .A2(n2668), .B1(n267), .B2(n901), .ZN(n1231) );
  NAND2_X2 U329 ( .A1(n627), .A2(n2395), .ZN(n1230) );
  NAND2_X2 U330 ( .A1(ready), .A2(i_start), .ZN(n627) );
  OAI22_X2 U331 ( .A1(n64), .A2(n913), .B1(n2335), .B2(n914), .ZN(n1229) );
  OAI22_X2 U332 ( .A1(n64), .A2(n915), .B1(n239), .B2(n914), .ZN(n1228) );
  OAI22_X2 U333 ( .A1(n2429), .A2(n539), .B1(n2427), .B2(n108), .ZN(n1227) );
  OAI22_X2 U334 ( .A1(n64), .A2(n916), .B1(n238), .B2(n914), .ZN(n1226) );
  OAI22_X2 U335 ( .A1(n64), .A2(n611), .B1(n241), .B2(n914), .ZN(n1225) );
  OAI22_X2 U336 ( .A1(n2424), .A2(n2669), .B1(n900), .B2(n719), .ZN(n1224) );
  OAI22_X2 U337 ( .A1(n2424), .A2(n2670), .B1(n719), .B2(n280), .ZN(n1223) );
  OAI22_X2 U338 ( .A1(n2424), .A2(n2671), .B1(n719), .B2(n278), .ZN(n1222) );
  OAI22_X2 U339 ( .A1(n2424), .A2(n2672), .B1(n719), .B2(n902), .ZN(n1221) );
  OAI22_X2 U340 ( .A1(n2424), .A2(n2673), .B1(n719), .B2(n903), .ZN(n1220) );
  OAI22_X2 U341 ( .A1(n2424), .A2(n2674), .B1(n719), .B2(n271), .ZN(n1219) );
  OAI22_X2 U342 ( .A1(n2424), .A2(n2675), .B1(n719), .B2(n270), .ZN(n1218) );
  OAI22_X2 U343 ( .A1(n2424), .A2(n2676), .B1(n2422), .B2(n904), .ZN(n1217) );
  OAI22_X2 U344 ( .A1(n2424), .A2(n2677), .B1(n719), .B2(n905), .ZN(n1216) );
  OAI22_X2 U345 ( .A1(n2424), .A2(n2678), .B1(n2422), .B2(n906), .ZN(n1215) );
  OAI22_X2 U346 ( .A1(n2424), .A2(n2679), .B1(n2422), .B2(n907), .ZN(n1214) );
  OAI22_X2 U347 ( .A1(n2424), .A2(n2680), .B1(n2422), .B2(n259), .ZN(n1213) );
  OAI22_X2 U348 ( .A1(n2424), .A2(n2681), .B1(n2422), .B2(n908), .ZN(n1212) );
  OAI22_X2 U349 ( .A1(n2424), .A2(n2682), .B1(n2422), .B2(n245), .ZN(n1211) );
  OAI22_X2 U350 ( .A1(n2424), .A2(n2683), .B1(n2422), .B2(n244), .ZN(n1210) );
  OAI22_X2 U351 ( .A1(n2425), .A2(n2684), .B1(n2422), .B2(n266), .ZN(n1209) );
  OAI22_X2 U352 ( .A1(n2425), .A2(n2685), .B1(n2422), .B2(n265), .ZN(n1208) );
  OAI22_X2 U353 ( .A1(n2425), .A2(n2686), .B1(n2422), .B2(n909), .ZN(n1207) );
  OAI22_X2 U354 ( .A1(n2425), .A2(n2687), .B1(n2422), .B2(n254), .ZN(n1206) );
  OAI22_X2 U355 ( .A1(n2425), .A2(n2688), .B1(n2422), .B2(n910), .ZN(n1205) );
  OAI22_X2 U356 ( .A1(n2425), .A2(n2689), .B1(n2422), .B2(n911), .ZN(n1204) );
  OAI22_X2 U357 ( .A1(n2423), .A2(n2690), .B1(n2422), .B2(n247), .ZN(n1203) );
  OAI22_X2 U358 ( .A1(n2424), .A2(n2691), .B1(n2422), .B2(n246), .ZN(n1202) );
  OAI22_X2 U359 ( .A1(n2423), .A2(n2692), .B1(n2422), .B2(n264), .ZN(n1201) );
  OAI22_X2 U360 ( .A1(n2423), .A2(n2693), .B1(n2422), .B2(n263), .ZN(n1200) );
  OAI22_X2 U361 ( .A1(n2423), .A2(n2694), .B1(n2422), .B2(n912), .ZN(n1199) );
  OAI22_X2 U362 ( .A1(n2424), .A2(n2695), .B1(n2422), .B2(n249), .ZN(n1198) );
  OAI22_X2 U363 ( .A1(n2424), .A2(n2696), .B1(n2422), .B2(n257), .ZN(n1197) );
  OAI22_X2 U364 ( .A1(n2424), .A2(n2697), .B1(n2422), .B2(n256), .ZN(n1196) );
  OAI22_X2 U365 ( .A1(n2424), .A2(n2698), .B1(n2422), .B2(n243), .ZN(n1195) );
  OAI22_X2 U366 ( .A1(n2424), .A2(n2699), .B1(n2422), .B2(n242), .ZN(n1194) );
  OAI22_X2 U367 ( .A1(n2424), .A2(n2700), .B1(n2422), .B2(n267), .ZN(n1193) );
  XOR2_X2 U368 ( .A(n933), .B(n940), .Z(n769) );
  XOR2_X2 U369 ( .A(reg_b[31]), .B(reg_a[31]), .Z(n940) );
  AOI22_X2 U374 ( .A1(n957), .A2(n958), .B1(n959), .B2(n960), .ZN(n942) );
  NAND2_X2 U376 ( .A1(n962), .A2(n958), .ZN(n953) );
  OAI22_X2 U377 ( .A1(n64), .A2(n963), .B1(n240), .B2(n914), .ZN(n1192) );
  OAI22_X2 U378 ( .A1(n64), .A2(n964), .B1(n105), .B2(n914), .ZN(n1191) );
  NAND4_X2 U379 ( .A1(n2394), .A2(n966), .A3(n967), .A4(n901), .ZN(n914) );
  NAND2_X2 U381 ( .A1(n2422), .A2(n613), .ZN(n977) );
  OAI22_X2 U383 ( .A1(n44), .A2(n969), .B1(n3116), .B2(n970), .ZN(n1190) );
  AOI22_X2 U384 ( .A1(n971), .A2(n972), .B1(n973), .B2(n974), .ZN(n969) );
  AOI22_X2 U386 ( .A1(n366), .A2(n2384), .B1(n367), .B2(n1114), .ZN(n971) );
  OAI211_X2 U387 ( .C1(n3117), .C2(n970), .A(n1115), .B(n1116), .ZN(n1189) );
  NAND4_X2 U388 ( .A1(n976), .A2(n1117), .A3(n2020), .A4(n1118), .ZN(n1115) );
  OAI211_X2 U389 ( .C1(n3118), .C2(n970), .A(n1119), .B(n1116), .ZN(n1188) );
  OAI22_X2 U392 ( .A1(n44), .A2(n974), .B1(n3119), .B2(n970), .ZN(n1187) );
  NAND2_X2 U393 ( .A1(n44), .A2(n2394), .ZN(n970) );
  NAND2_X2 U394 ( .A1(n68), .A2(n2434), .ZN(n1118) );
  OAI221_X2 U395 ( .B1(n2412), .B2(n580), .C1(n298), .C2(n2407), .A(n1121), 
        .ZN(n1186) );
  OAI221_X2 U398 ( .B1(n2412), .B2(n579), .C1(n345), .C2(n2407), .A(n1122), 
        .ZN(n1185) );
  OAI221_X2 U401 ( .B1(n2412), .B2(n578), .C1(n390), .C2(n2407), .A(n1298), 
        .ZN(n1184) );
  OAI22_X2 U403 ( .A1(n1300), .A2(n2382), .B1(n1295), .B2(n2378), .ZN(n615) );
  AOI22_X2 U404 ( .A1(n2387), .A2(sdata[1]), .B1(n2377), .B2(sdata[0]), .ZN(
        n1295) );
  OAI221_X2 U405 ( .B1(n2412), .B2(n577), .C1(n387), .C2(n2407), .A(n1303), 
        .ZN(n1183) );
  OAI221_X2 U408 ( .B1(n2412), .B2(n576), .C1(n386), .C2(n2407), .A(n1305), 
        .ZN(n1182) );
  OAI22_X2 U410 ( .A1(n296), .A2(n2374), .B1(n297), .B2(n2370), .ZN(n620) );
  OAI22_X2 U411 ( .A1(n1308), .A2(n2382), .B1(n2379), .B2(n1300), .ZN(n1307)
         );
  AOI22_X2 U412 ( .A1(n2387), .A2(sdata[2]), .B1(n2377), .B2(sdata[1]), .ZN(
        n1300) );
  OAI221_X2 U413 ( .B1(n2412), .B2(n575), .C1(n385), .C2(n2407), .A(n1309), 
        .ZN(n1181) );
  NOR4_X2 U415 ( .A1(n294), .A2(n2341), .A3(n361), .A4(n2343), .ZN(n622) );
  OAI221_X2 U416 ( .B1(n2412), .B2(n574), .C1(n388), .C2(n2407), .A(n1312), 
        .ZN(n1180) );
  XNOR2_X2 U418 ( .A(n1313), .B(n1314), .ZN(n917) );
  AOI22_X2 U421 ( .A1(n294), .A2(n2341), .B1(n1320), .B2(n293), .ZN(n1319) );
  OAI221_X2 U422 ( .B1(n2412), .B2(n573), .C1(n389), .C2(n2407), .A(n1321), 
        .ZN(n1179) );
  XNOR2_X2 U424 ( .A(n1322), .B(n1323), .ZN(n904) );
  OAI211_X2 U425 ( .C1(n2021), .C2(n1324), .A(n1318), .B(n1325), .ZN(n724) );
  AOI22_X2 U426 ( .A1(n293), .A2(n2341), .B1(n343), .B2(n1320), .ZN(n1325) );
  OAI221_X2 U427 ( .B1(n2412), .B2(n572), .C1(n391), .C2(n2407), .A(n1326), 
        .ZN(n1178) );
  XOR2_X2 U429 ( .A(n1327), .B(n1328), .Z(n905) );
  OAI221_X2 U431 ( .B1(n1330), .B2(n1331), .C1(n2342), .C2(n1332), .A(n1333), 
        .ZN(n725) );
  AOI22_X2 U432 ( .A1(n294), .A2(n361), .B1(n293), .B2(n2343), .ZN(n1333) );
  OAI22_X2 U433 ( .A1(n295), .A2(n2374), .B1(n296), .B2(n2372), .ZN(n1324) );
  OAI22_X2 U434 ( .A1(n1335), .A2(n2382), .B1(n2378), .B2(n1308), .ZN(n1334)
         );
  OAI221_X2 U435 ( .B1(n2411), .B2(n571), .C1(n392), .C2(n2407), .A(n1336), 
        .ZN(n1177) );
  XNOR2_X2 U437 ( .A(n1337), .B(n1338), .ZN(n906) );
  OAI221_X2 U438 ( .B1(n1330), .B2(n1332), .C1(n2342), .C2(n1339), .A(n1340), 
        .ZN(n726) );
  AOI22_X2 U439 ( .A1(n293), .A2(n361), .B1(n343), .B2(n2343), .ZN(n1340) );
  OAI22_X2 U440 ( .A1(n344), .A2(n2374), .B1(n295), .B2(n2372), .ZN(n1341) );
  OAI221_X2 U441 ( .B1(n2411), .B2(n570), .C1(n342), .C2(n2408), .A(n1342), 
        .ZN(n1176) );
  XOR2_X2 U443 ( .A(n1343), .B(n1344), .Z(n907) );
  OAI221_X2 U445 ( .B1(n1330), .B2(n1339), .C1(n2342), .C2(n1346), .A(n1347), 
        .ZN(n727) );
  AOI22_X2 U446 ( .A1(n343), .A2(n361), .B1(n356), .B2(n2343), .ZN(n1347) );
  OAI22_X2 U447 ( .A1(n358), .A2(n2374), .B1(n344), .B2(n2372), .ZN(n1331) );
  OAI221_X2 U448 ( .B1(n2411), .B2(n569), .C1(n322), .C2(n2408), .A(n1348), 
        .ZN(n1175) );
  XOR2_X2 U450 ( .A(n1349), .B(n1350), .Z(n918) );
  OAI221_X2 U451 ( .B1(n1330), .B2(n1346), .C1(n2342), .C2(n1351), .A(n1352), 
        .ZN(n728) );
  AOI22_X2 U452 ( .A1(n356), .A2(n361), .B1(n287), .B2(n2343), .ZN(n1352) );
  OAI22_X2 U453 ( .A1(n357), .A2(n2374), .B1(n358), .B2(n2371), .ZN(n1332) );
  OAI221_X2 U454 ( .B1(n2411), .B2(n568), .C1(n339), .C2(n2408), .A(n1353), 
        .ZN(n1174) );
  XOR2_X2 U456 ( .A(n1354), .B(n1355), .Z(n908) );
  OAI221_X2 U458 ( .B1(n1330), .B2(n1351), .C1(n2342), .C2(n1357), .A(n1358), 
        .ZN(n729) );
  AOI22_X2 U459 ( .A1(n287), .A2(n361), .B1(n340), .B2(n2343), .ZN(n1358) );
  OAI222_X2 U460 ( .A1(n357), .A2(n2370), .B1(n295), .B2(n2383), .C1(n355), 
        .C2(n2373), .ZN(n1339) );
  OAI222_X2 U461 ( .A1(n2378), .A2(n1335), .B1(n1308), .B2(n2439), .C1(n1360), 
        .C2(n2381), .ZN(n1359) );
  OAI221_X2 U463 ( .B1(n2411), .B2(n567), .C1(n338), .C2(n2408), .A(n1361), 
        .ZN(n1173) );
  XOR2_X2 U465 ( .A(n494), .B(n1362), .Z(n919) );
  OAI221_X2 U466 ( .B1(n1330), .B2(n1357), .C1(n2342), .C2(n1363), .A(n1364), 
        .ZN(n730) );
  AOI22_X2 U467 ( .A1(n340), .A2(n361), .B1(n312), .B2(n2343), .ZN(n1364) );
  OAI222_X2 U468 ( .A1(n355), .A2(n2370), .B1(n344), .B2(n2383), .C1(n341), 
        .C2(n2373), .ZN(n1346) );
  OAI222_X2 U469 ( .A1(n2378), .A2(n1360), .B1(n1335), .B2(n2439), .C1(n1366), 
        .C2(n2381), .ZN(n1365) );
  OAI221_X2 U471 ( .B1(n2411), .B2(n566), .C1(n337), .C2(n2408), .A(n1367), 
        .ZN(n1172) );
  XOR2_X2 U473 ( .A(n1368), .B(n1369), .Z(n920) );
  OAI221_X2 U475 ( .B1(n1330), .B2(n1363), .C1(n2342), .C2(n1371), .A(n1372), 
        .ZN(n731) );
  AOI22_X2 U476 ( .A1(n312), .A2(n361), .B1(n309), .B2(n2343), .ZN(n1372) );
  OAI222_X2 U477 ( .A1(n341), .A2(n2370), .B1(n358), .B2(n2383), .C1(n313), 
        .C2(n2373), .ZN(n1351) );
  OAI222_X2 U478 ( .A1(n2378), .A2(n1366), .B1(n1360), .B2(n2439), .C1(n1374), 
        .C2(n2381), .ZN(n1373) );
  OAI221_X2 U480 ( .B1(n2411), .B2(n565), .C1(n336), .C2(n2408), .A(n1375), 
        .ZN(n1171) );
  XOR2_X2 U482 ( .A(n955), .B(n1376), .Z(n921) );
  OAI221_X2 U483 ( .B1(n1330), .B2(n1371), .C1(n2342), .C2(n1377), .A(n1378), 
        .ZN(n732) );
  AOI22_X2 U484 ( .A1(n309), .A2(n361), .B1(n306), .B2(n2343), .ZN(n1378) );
  OAI222_X2 U485 ( .A1(n313), .A2(n2370), .B1(n357), .B2(n2383), .C1(n310), 
        .C2(n2373), .ZN(n1357) );
  OAI222_X2 U486 ( .A1(n2379), .A2(n1374), .B1(n1366), .B2(n2439), .C1(n1380), 
        .C2(n2381), .ZN(n1379) );
  OAI221_X2 U488 ( .B1(n2411), .B2(n564), .C1(n335), .C2(n2408), .A(n1381), 
        .ZN(n1170) );
  XNOR2_X2 U490 ( .A(n1382), .B(n1383), .ZN(n922) );
  NAND2_X2 U492 ( .A1(n1385), .A2(n1386), .ZN(n955) );
  OAI221_X2 U493 ( .B1(n1330), .B2(n1377), .C1(n2342), .C2(n1387), .A(n1388), 
        .ZN(n733) );
  AOI22_X2 U494 ( .A1(n306), .A2(n361), .B1(n303), .B2(n2343), .ZN(n1388) );
  OAI222_X2 U495 ( .A1(n310), .A2(n2370), .B1(n355), .B2(n2383), .C1(n308), 
        .C2(n2373), .ZN(n1363) );
  OAI222_X2 U496 ( .A1(n2378), .A2(n1380), .B1(n1374), .B2(n2439), .C1(n1390), 
        .C2(n2381), .ZN(n1389) );
  OAI221_X2 U498 ( .B1(n2411), .B2(n563), .C1(n380), .C2(n2408), .A(n1391), 
        .ZN(n1169) );
  XOR2_X2 U500 ( .A(n1392), .B(n1393), .Z(n909) );
  OAI221_X2 U501 ( .B1(n1330), .B2(n1387), .C1(n2342), .C2(n1394), .A(n1395), 
        .ZN(n734) );
  AOI22_X2 U502 ( .A1(n303), .A2(n361), .B1(n311), .B2(n2343), .ZN(n1395) );
  OAI222_X2 U503 ( .A1(n308), .A2(n2370), .B1(n341), .B2(n2383), .C1(n316), 
        .C2(n2373), .ZN(n1371) );
  OAI222_X2 U504 ( .A1(n2378), .A2(n1390), .B1(n1380), .B2(n2439), .C1(n1397), 
        .C2(n2381), .ZN(n1396) );
  OAI221_X2 U506 ( .B1(n2411), .B2(n562), .C1(n381), .C2(n2408), .A(n1398), 
        .ZN(n1168) );
  XOR2_X2 U508 ( .A(n1399), .B(n1400), .Z(n923) );
  AOI221_X2 U510 ( .B1(n1402), .B2(n1403), .C1(n1403), .C2(n1404), .A(n1405), 
        .ZN(n1392) );
  AOI221_X2 U511 ( .B1(n2341), .B2(n300), .C1(n1320), .C2(n315), .A(n1406), 
        .ZN(n736) );
  OAI22_X2 U512 ( .A1(n1377), .A2(n1318), .B1(n1387), .B2(n2021), .ZN(n1406)
         );
  OAI222_X2 U513 ( .A1(n316), .A2(n2371), .B1(n313), .B2(n2383), .C1(n321), 
        .C2(n2373), .ZN(n1377) );
  OAI222_X2 U514 ( .A1(n2378), .A2(n1397), .B1(n1390), .B2(n2439), .C1(n1408), 
        .C2(n2381), .ZN(n1407) );
  OAI221_X2 U516 ( .B1(n2411), .B2(n561), .C1(n379), .C2(n2408), .A(n1409), 
        .ZN(n1167) );
  XNOR2_X2 U518 ( .A(n1410), .B(n1411), .ZN(n910) );
  AOI221_X2 U519 ( .B1(n2341), .B2(n315), .C1(n1320), .C2(n320), .A(n1412), 
        .ZN(n737) );
  OAI22_X2 U520 ( .A1(n1387), .A2(n1318), .B1(n1394), .B2(n2021), .ZN(n1412)
         );
  OAI222_X2 U521 ( .A1(n321), .A2(n2371), .B1(n310), .B2(n2383), .C1(n319), 
        .C2(n2373), .ZN(n1387) );
  OAI222_X2 U522 ( .A1(n2378), .A2(n1408), .B1(n1397), .B2(n2439), .C1(n1414), 
        .C2(n2381), .ZN(n1413) );
  OAI221_X2 U524 ( .B1(n2410), .B2(n560), .C1(n378), .C2(n2408), .A(n1416), 
        .ZN(n1166) );
  XOR2_X2 U526 ( .A(n1417), .B(n1418), .Z(n911) );
  OAI221_X2 U528 ( .B1(n1420), .B2(n1421), .C1(n1421), .C2(n1422), .A(n1423), 
        .ZN(n1410) );
  NAND2_X2 U529 ( .A1(n1424), .A2(n1425), .ZN(n1421) );
  AOI221_X2 U530 ( .B1(n2341), .B2(n320), .C1(n1320), .C2(n318), .A(n1426), 
        .ZN(n739) );
  OAI22_X2 U531 ( .A1(n1394), .A2(n1318), .B1(n1415), .B2(n2021), .ZN(n1426)
         );
  OAI222_X2 U532 ( .A1(n319), .A2(n2371), .B1(n308), .B2(n2383), .C1(n327), 
        .C2(n2373), .ZN(n1394) );
  OAI222_X2 U533 ( .A1(n2378), .A2(n1414), .B1(n1408), .B2(n2439), .C1(n1428), 
        .C2(n2381), .ZN(n1427) );
  OAI221_X2 U535 ( .B1(n2410), .B2(n559), .C1(n377), .C2(n2409), .A(n1430), 
        .ZN(n1165) );
  XOR2_X2 U537 ( .A(n1431), .B(n1432), .Z(n924) );
  AOI221_X2 U538 ( .B1(n2341), .B2(n318), .C1(n1320), .C2(n326), .A(n1433), 
        .ZN(n740) );
  OAI22_X2 U539 ( .A1(n1415), .A2(n1318), .B1(n1429), .B2(n2021), .ZN(n1433)
         );
  OAI222_X2 U540 ( .A1(n327), .A2(n2371), .B1(n316), .B2(n2383), .C1(n325), 
        .C2(n2373), .ZN(n1415) );
  OAI222_X2 U541 ( .A1(n2378), .A2(n1428), .B1(n1414), .B2(n2439), .C1(n1435), 
        .C2(n2381), .ZN(n1434) );
  OAI221_X2 U543 ( .B1(n2410), .B2(n558), .C1(n376), .C2(n2409), .A(n1437), 
        .ZN(n1164) );
  XNOR2_X2 U545 ( .A(n1438), .B(n1439), .ZN(n925) );
  OAI211_X2 U547 ( .C1(n248), .C2(n1441), .A(n1442), .B(n495), .ZN(n1431) );
  AOI221_X2 U549 ( .B1(n2341), .B2(n326), .C1(n1320), .C2(n324), .A(n1446), 
        .ZN(n742) );
  OAI22_X2 U550 ( .A1(n1429), .A2(n1318), .B1(n1436), .B2(n2021), .ZN(n1446)
         );
  OAI222_X2 U551 ( .A1(n325), .A2(n2371), .B1(n321), .B2(n2383), .C1(n329), 
        .C2(n2373), .ZN(n1429) );
  OAI222_X2 U552 ( .A1(n2378), .A2(n1435), .B1(n1428), .B2(n2439), .C1(n1448), 
        .C2(n2381), .ZN(n1447) );
  OAI221_X2 U554 ( .B1(n2410), .B2(n557), .C1(n375), .C2(n2409), .A(n1450), 
        .ZN(n1163) );
  XOR2_X2 U556 ( .A(n1451), .B(n1452), .Z(n926) );
  AOI221_X2 U557 ( .B1(n2341), .B2(n324), .C1(n1320), .C2(n328), .A(n1453), 
        .ZN(n743) );
  OAI22_X2 U558 ( .A1(n1436), .A2(n1318), .B1(n1449), .B2(n2021), .ZN(n1453)
         );
  OAI222_X2 U559 ( .A1(n329), .A2(n2371), .B1(n319), .B2(n2383), .C1(n334), 
        .C2(n2373), .ZN(n1436) );
  OAI222_X2 U560 ( .A1(n2378), .A2(n1448), .B1(n1435), .B2(n2440), .C1(n1455), 
        .C2(n2381), .ZN(n1454) );
  OAI221_X2 U562 ( .B1(n2410), .B2(n556), .C1(n374), .C2(n2409), .A(n1457), 
        .ZN(n1162) );
  XNOR2_X2 U564 ( .A(n1458), .B(n1459), .ZN(n927) );
  OAI221_X2 U566 ( .B1(n1385), .B2(n1461), .C1(n1461), .C2(n1386), .A(n954), 
        .ZN(n1451) );
  NAND2_X2 U569 ( .A1(n1466), .A2(n1467), .ZN(n1322) );
  AOI221_X2 U572 ( .B1(n2341), .B2(n328), .C1(n1472), .C2(n1320), .A(n1473), 
        .ZN(n745) );
  OAI22_X2 U573 ( .A1(n1449), .A2(n1318), .B1(n1456), .B2(n2021), .ZN(n1473)
         );
  OAI222_X2 U574 ( .A1(n334), .A2(n2370), .B1(n327), .B2(n2383), .C1(n333), 
        .C2(n2373), .ZN(n1449) );
  OAI222_X2 U575 ( .A1(n2379), .A2(n1455), .B1(n1448), .B2(n2440), .C1(n1475), 
        .C2(n2381), .ZN(n1474) );
  OAI221_X2 U577 ( .B1(n2410), .B2(n555), .C1(n373), .C2(n2409), .A(n1477), 
        .ZN(n1161) );
  XOR2_X2 U579 ( .A(n1478), .B(n1479), .Z(n912) );
  AOI221_X2 U580 ( .B1(n1472), .B2(n2341), .C1(n1480), .C2(n1320), .A(n1481), 
        .ZN(n746) );
  OAI22_X2 U581 ( .A1(n1456), .A2(n1318), .B1(n1482), .B2(n2021), .ZN(n1481)
         );
  OAI222_X2 U582 ( .A1(n333), .A2(n2370), .B1(n325), .B2(n2383), .C1(n354), 
        .C2(n2374), .ZN(n1456) );
  OAI222_X2 U583 ( .A1(n2379), .A2(n1475), .B1(n1455), .B2(n2440), .C1(n1484), 
        .C2(n2382), .ZN(n1483) );
  OAI221_X2 U585 ( .B1(n2410), .B2(n554), .C1(n372), .C2(n2409), .A(n1486), 
        .ZN(n1160) );
  XNOR2_X2 U587 ( .A(n1487), .B(n1488), .ZN(n928) );
  OAI211_X2 U589 ( .C1(n1490), .C2(n1491), .A(n1492), .B(n1493), .ZN(n1478) );
  OR2_X2 U594 ( .A1(n1402), .A2(n1404), .ZN(n1337) );
  AND4_X2 U595 ( .A1(n272), .A2(n1469), .A3(n1499), .A4(n1500), .ZN(n1404) );
  AOI221_X2 U599 ( .B1(n361), .B2(n328), .C1(n1472), .C2(n2343), .A(n332), 
        .ZN(n748) );
  AOI22_X2 U600 ( .A1(n2341), .A2(n1480), .B1(n1320), .B2(n1508), .ZN(n1507)
         );
  OAI222_X2 U601 ( .A1(n354), .A2(n2370), .B1(n329), .B2(n2383), .C1(n353), 
        .C2(n2374), .ZN(n1482) );
  OAI222_X2 U602 ( .A1(n2379), .A2(n1484), .B1(n1475), .B2(n2440), .C1(n1511), 
        .C2(n2382), .ZN(n1510) );
  OAI221_X2 U604 ( .B1(n2410), .B2(n553), .C1(n370), .C2(n2409), .A(n1513), 
        .ZN(n1159) );
  XOR2_X2 U606 ( .A(n1514), .B(n1515), .Z(n929) );
  AOI221_X2 U607 ( .B1(n1508), .B2(n2341), .C1(n1516), .C2(n1320), .A(n331), 
        .ZN(n750) );
  AOI22_X2 U608 ( .A1(n361), .A2(n1472), .B1(n2343), .B2(n1480), .ZN(n1517) );
  OAI222_X2 U609 ( .A1(n2371), .A2(n1509), .B1(n2383), .B2(n1476), .C1(n2374), 
        .C2(n1518), .ZN(n1472) );
  OAI222_X2 U610 ( .A1(n2379), .A2(n1511), .B1(n1484), .B2(n2440), .C1(n1519), 
        .C2(n2382), .ZN(n1476) );
  OAI221_X2 U612 ( .B1(n2410), .B2(n552), .C1(n535), .C2(n2409), .A(n1520), 
        .ZN(n1158) );
  XNOR2_X2 U614 ( .A(n1521), .B(n1522), .ZN(n930) );
  AND3_X2 U616 ( .A1(n961), .A2(n1524), .A3(n1525), .ZN(n1514) );
  AOI22_X2 U617 ( .A1(n1526), .A2(n1463), .B1(n521), .B2(n1464), .ZN(n1525) );
  NAND2_X2 U618 ( .A1(n1527), .A2(n1528), .ZN(n1464) );
  NAND2_X2 U622 ( .A1(n1530), .A2(n1531), .ZN(n1462) );
  NAND2_X2 U624 ( .A1(n496), .A2(n1533), .ZN(n1471) );
  OR3_X2 U625 ( .A1(n498), .A2(n1534), .A3(n494), .ZN(n1533) );
  NAND4_X2 U626 ( .A1(n501), .A2(n521), .A3(n1425), .A4(n1349), .ZN(n1524) );
  NAND2_X2 U627 ( .A1(n1420), .A2(n1422), .ZN(n1349) );
  NAND4_X2 U628 ( .A1(n1465), .A2(n1469), .A3(n1468), .A4(n277), .ZN(n1422) );
  NAND2_X2 U630 ( .A1(n1536), .A2(n1537), .ZN(n1470) );
  AND4_X2 U632 ( .A1(n1323), .A2(n1328), .A3(n1338), .A4(n1344), .ZN(n1465) );
  NOR4_X2 U634 ( .A1(n482), .A2(n490), .A3(n494), .A4(n498), .ZN(n1425) );
  NAND2_X2 U636 ( .A1(n1424), .A2(n1463), .ZN(n1461) );
  AND4_X2 U637 ( .A1(n1438), .A2(n1432), .A3(n1418), .A4(n1411), .ZN(n1463) );
  AND4_X2 U638 ( .A1(n1400), .A2(n1393), .A3(n1382), .A4(n1376), .ZN(n1424) );
  OAI221_X2 U640 ( .B1(n350), .B2(n1330), .C1(n349), .C2(n2342), .A(n1545), 
        .ZN(n751) );
  AOI22_X2 U641 ( .A1(n361), .A2(n1480), .B1(n2343), .B2(n1508), .ZN(n1545) );
  OAI222_X2 U642 ( .A1(n2371), .A2(n1518), .B1(n2383), .B2(n1485), .C1(n2374), 
        .C2(n1546), .ZN(n1480) );
  OAI222_X2 U643 ( .A1(n2379), .A2(n1519), .B1(n1511), .B2(n2440), .C1(n1547), 
        .C2(n2382), .ZN(n1485) );
  OAI221_X2 U645 ( .B1(n2410), .B2(n551), .C1(n384), .C2(n2409), .A(n1548), 
        .ZN(n1157) );
  XOR2_X2 U647 ( .A(n962), .B(n1549), .Z(n931) );
  OAI221_X2 U648 ( .B1(n349), .B2(n1330), .C1(n348), .C2(n2342), .A(n1550), 
        .ZN(n752) );
  AOI22_X2 U649 ( .A1(n361), .A2(n1508), .B1(n2343), .B2(n1516), .ZN(n1550) );
  OAI222_X2 U651 ( .A1(n2371), .A2(n1546), .B1(n2383), .B2(n1512), .C1(n2374), 
        .C2(n1553), .ZN(n1508) );
  OAI222_X2 U652 ( .A1(n2379), .A2(n1547), .B1(n1519), .B2(n2440), .C1(n1554), 
        .C2(n2382), .ZN(n1512) );
  OAI221_X2 U655 ( .B1(n2410), .B2(n550), .C1(n534), .C2(n2409), .A(n1556), 
        .ZN(n1156) );
  XNOR2_X2 U658 ( .A(n1557), .B(n958), .ZN(n932) );
  XNOR2_X2 U659 ( .A(reg_a[30]), .B(n538), .ZN(n958) );
  AND2_X2 U661 ( .A1(reg_b[29]), .A2(reg_a[29]), .ZN(n957) );
  XOR2_X2 U662 ( .A(reg_a[29]), .B(reg_b[29]), .Z(n962) );
  OAI211_X2 U663 ( .C1(n495), .C2(n1558), .A(n527), .B(n1559), .ZN(n1549) );
  NAND2_X2 U665 ( .A1(n1544), .A2(n1561), .ZN(n1495) );
  AOI22_X2 U667 ( .A1(reg_b[22]), .A2(reg_a[22]), .B1(n1438), .B2(n1440), .ZN(
        n1527) );
  AND2_X2 U668 ( .A1(reg_a[21]), .A2(reg_b[21]), .ZN(n1440) );
  AOI22_X2 U669 ( .A1(reg_b[24]), .A2(reg_a[24]), .B1(n1458), .B2(n1460), .ZN(
        n1544) );
  AND2_X2 U670 ( .A1(reg_b[23]), .A2(reg_a[23]), .ZN(n1460) );
  OR2_X2 U671 ( .A1(n1444), .A2(n1497), .ZN(n1441) );
  NAND4_X2 U672 ( .A1(n1382), .A2(n1376), .A3(n1541), .A4(n1369), .ZN(n1497)
         );
  XOR2_X2 U673 ( .A(reg_a[13]), .B(reg_b[13]), .Z(n1541) );
  AND2_X2 U676 ( .A1(n1534), .A2(n1562), .ZN(n1496) );
  OR3_X2 U677 ( .A1(n490), .A2(n1536), .A3(n482), .ZN(n1562) );
  AOI22_X2 U678 ( .A1(reg_b[10]), .A2(reg_a[10]), .B1(n1344), .B2(n1345), .ZN(
        n1536) );
  AND2_X2 U679 ( .A1(reg_b[9]), .A2(reg_a[9]), .ZN(n1345) );
  AOI22_X2 U680 ( .A1(reg_b[12]), .A2(reg_a[12]), .B1(n1355), .B2(n1356), .ZN(
        n1534) );
  AND2_X2 U681 ( .A1(reg_b[11]), .A2(reg_a[11]), .ZN(n1356) );
  AND2_X2 U682 ( .A1(n1538), .A2(n1563), .ZN(n1505) );
  OAI22_X2 U684 ( .A1(n487), .A2(n497), .B1(n1314), .B2(n1317), .ZN(n1540) );
  NAND2_X2 U685 ( .A1(reg_b[5]), .A2(reg_a[5]), .ZN(n1317) );
  AOI22_X2 U686 ( .A1(reg_b[8]), .A2(reg_a[8]), .B1(n1328), .B2(n1329), .ZN(
        n1538) );
  AND2_X2 U687 ( .A1(reg_b[7]), .A2(reg_a[7]), .ZN(n1329) );
  XOR2_X2 U691 ( .A(reg_a[6]), .B(n487), .Z(n1314) );
  XOR2_X2 U692 ( .A(reg_a[8]), .B(reg_b[8]), .Z(n1328) );
  XOR2_X2 U693 ( .A(reg_a[7]), .B(reg_b[7]), .Z(n1323) );
  NAND4_X2 U694 ( .A1(n1338), .A2(n1344), .A3(n1350), .A4(n1355), .ZN(n1506)
         );
  XOR2_X2 U695 ( .A(reg_a[12]), .B(reg_b[12]), .Z(n1355) );
  XOR2_X2 U696 ( .A(reg_a[11]), .B(reg_b[11]), .Z(n1350) );
  XOR2_X2 U697 ( .A(reg_a[10]), .B(reg_b[10]), .Z(n1344) );
  XOR2_X2 U698 ( .A(reg_a[9]), .B(reg_b[9]), .Z(n1338) );
  OAI22_X2 U699 ( .A1(n525), .A2(n526), .B1(n1488), .B2(n1489), .ZN(n1543) );
  NAND2_X2 U700 ( .A1(reg_b[25]), .A2(reg_a[25]), .ZN(n1489) );
  OAI22_X2 U701 ( .A1(n531), .A2(n536), .B1(n1522), .B2(n1523), .ZN(n952) );
  NAND2_X2 U702 ( .A1(reg_a[27]), .A2(reg_b[27]), .ZN(n1523) );
  OR3_X2 U703 ( .A1(n528), .A2(n523), .A3(n1491), .ZN(n1558) );
  NAND4_X2 U704 ( .A1(n1438), .A2(n1432), .A3(n1458), .A4(n1452), .ZN(n1491)
         );
  XOR2_X2 U705 ( .A(reg_a[23]), .B(reg_b[23]), .Z(n1452) );
  XOR2_X2 U706 ( .A(reg_a[24]), .B(reg_b[24]), .Z(n1458) );
  XNOR2_X2 U707 ( .A(reg_a[21]), .B(n517), .ZN(n1432) );
  XOR2_X2 U708 ( .A(reg_a[22]), .B(reg_b[22]), .Z(n1438) );
  XOR2_X2 U710 ( .A(reg_a[26]), .B(n525), .Z(n1488) );
  XOR2_X2 U711 ( .A(reg_a[25]), .B(n524), .Z(n1479) );
  XOR2_X2 U713 ( .A(reg_a[28]), .B(n531), .Z(n1522) );
  XOR2_X2 U714 ( .A(reg_a[27]), .B(n529), .Z(n1515) );
  AND2_X2 U716 ( .A1(n1529), .A2(n1565), .ZN(n1490) );
  AOI22_X2 U718 ( .A1(reg_b[18]), .A2(reg_a[18]), .B1(n1400), .B2(n507), .ZN(
        n1530) );
  NAND2_X2 U719 ( .A1(reg_a[17]), .A2(reg_b[17]), .ZN(n1401) );
  AOI22_X2 U720 ( .A1(reg_b[20]), .A2(reg_a[20]), .B1(n1418), .B2(n1419), .ZN(
        n1529) );
  AND2_X2 U721 ( .A1(reg_a[19]), .A2(reg_b[19]), .ZN(n1419) );
  NAND4_X2 U722 ( .A1(n1418), .A2(n1411), .A3(n1400), .A4(n1393), .ZN(n1444)
         );
  XOR2_X2 U723 ( .A(reg_a[17]), .B(reg_b[17]), .Z(n1393) );
  XOR2_X2 U724 ( .A(reg_a[18]), .B(reg_b[18]), .Z(n1400) );
  XOR2_X2 U725 ( .A(reg_a[19]), .B(reg_b[19]), .Z(n1411) );
  XOR2_X2 U726 ( .A(reg_a[20]), .B(reg_b[20]), .Z(n1418) );
  AND2_X2 U727 ( .A1(n1532), .A2(n1566), .ZN(n1498) );
  OAI22_X2 U729 ( .A1(n499), .A2(n500), .B1(n498), .B2(n1370), .ZN(n1535) );
  NAND2_X2 U730 ( .A1(reg_b[13]), .A2(reg_a[13]), .ZN(n1370) );
  XOR2_X2 U731 ( .A(reg_a[14]), .B(reg_b[14]), .Z(n1369) );
  XNOR2_X2 U732 ( .A(reg_a[15]), .B(n502), .ZN(n1376) );
  AOI22_X2 U733 ( .A1(reg_b[16]), .A2(reg_a[16]), .B1(n1382), .B2(n1384), .ZN(
        n1532) );
  AND2_X2 U734 ( .A1(reg_a[15]), .A2(reg_b[15]), .ZN(n1384) );
  XOR2_X2 U735 ( .A(reg_a[16]), .B(reg_b[16]), .Z(n1382) );
  OAI222_X2 U736 ( .A1(n348), .A2(n1330), .B1(n350), .B2(n1318), .C1(n1567), 
        .C2(n1551), .ZN(n753) );
  AOI22_X2 U737 ( .A1(n1552), .A2(n1568), .B1(n364), .B2(n1555), .ZN(n1567) );
  OAI222_X2 U738 ( .A1(n2371), .A2(n1569), .B1(n2383), .B2(n1518), .C1(n1570), 
        .C2(n2374), .ZN(n1555) );
  OAI222_X2 U739 ( .A1(n2379), .A2(n1571), .B1(n1554), .B2(n2440), .C1(n1572), 
        .C2(n2382), .ZN(n1518) );
  OAI222_X2 U740 ( .A1(n1573), .A2(n2370), .B1(n2383), .B2(n1553), .C1(n1574), 
        .C2(n2374), .ZN(n1568) );
  OAI222_X2 U744 ( .A1(n2371), .A2(n1553), .B1(n2383), .B2(n1509), .C1(n2374), 
        .C2(n1569), .ZN(n1516) );
  OAI222_X2 U745 ( .A1(n2379), .A2(n1577), .B1(n1578), .B2(n2440), .C1(n2382), 
        .C2(n351), .ZN(n1569) );
  OAI222_X2 U746 ( .A1(n2379), .A2(n1554), .B1(n1547), .B2(n2440), .C1(n1571), 
        .C2(n2382), .ZN(n1509) );
  OAI222_X2 U749 ( .A1(n2379), .A2(n1578), .B1(n1572), .B2(n2440), .C1(n1577), 
        .C2(n2382), .ZN(n1553) );
  NAND2_X2 U750 ( .A1(n1552), .A2(n1551), .ZN(n1330) );
  NAND2_X2 U753 ( .A1(n973), .A2(n2384), .ZN(n1552) );
  OAI222_X2 U754 ( .A1(n1570), .A2(n2370), .B1(n2384), .B2(n1546), .C1(n1573), 
        .C2(n2373), .ZN(n1580) );
  OAI222_X2 U758 ( .A1(n2378), .A2(n1572), .B1(n1571), .B2(n2439), .C1(n1578), 
        .C2(n2381), .ZN(n1546) );
  NAND2_X2 U763 ( .A1(n1583), .A2(n973), .ZN(n974) );
  AND2_X2 U764 ( .A1(n1584), .A2(n366), .ZN(n973) );
  NAND2_X2 U765 ( .A1(n1585), .A2(n1575), .ZN(n1120) );
  XOR2_X2 U766 ( .A(n373), .B(n2019), .Z(n1585) );
  XOR2_X2 U767 ( .A(n374), .B(n2019), .Z(n1584) );
  XOR2_X2 U768 ( .A(n375), .B(n2019), .Z(n1583) );
  XOR2_X2 U776 ( .A(n372), .B(n2334), .Z(n1114) );
  NAND2_X2 U777 ( .A1(n1587), .A2(n2438), .ZN(n1117) );
  XOR2_X2 U778 ( .A(n370), .B(n2019), .Z(n1587) );
  NAND2_X2 U780 ( .A1(n2377), .A2(n976), .ZN(n1301) );
  XOR2_X2 U783 ( .A(n535), .B(n2019), .Z(n1589) );
  XOR2_X2 U784 ( .A(n384), .B(n2019), .Z(n976) );
  OAI22_X2 U789 ( .A1(n298), .A2(n966), .B1(n2390), .B2(n118), .ZN(n1155) );
  OAI22_X2 U790 ( .A1(n345), .A2(n966), .B1(n2390), .B2(n117), .ZN(n1154) );
  OAI22_X2 U791 ( .A1(n390), .A2(n966), .B1(n2390), .B2(n116), .ZN(n1153) );
  OAI22_X2 U792 ( .A1(n387), .A2(n966), .B1(n2390), .B2(n115), .ZN(n1152) );
  OAI22_X2 U793 ( .A1(n386), .A2(n966), .B1(n2390), .B2(n114), .ZN(n1151) );
  OAI22_X2 U794 ( .A1(n385), .A2(n966), .B1(n2390), .B2(n113), .ZN(n1150) );
  OAI22_X2 U795 ( .A1(n388), .A2(n966), .B1(n2390), .B2(n112), .ZN(n1149) );
  OAI22_X2 U796 ( .A1(n389), .A2(n2389), .B1(n2390), .B2(n111), .ZN(n1148) );
  OAI22_X2 U797 ( .A1(n391), .A2(n2389), .B1(n2390), .B2(n143), .ZN(n1147) );
  OAI22_X2 U798 ( .A1(n392), .A2(n2389), .B1(n2390), .B2(n142), .ZN(n1146) );
  OAI22_X2 U799 ( .A1(n342), .A2(n2389), .B1(n2390), .B2(n141), .ZN(n1145) );
  OAI22_X2 U800 ( .A1(n322), .A2(n2388), .B1(n2390), .B2(n140), .ZN(n1144) );
  OAI22_X2 U801 ( .A1(n339), .A2(n2388), .B1(n2390), .B2(n139), .ZN(n1143) );
  OAI22_X2 U802 ( .A1(n338), .A2(n2388), .B1(n2390), .B2(n138), .ZN(n1142) );
  OAI22_X2 U803 ( .A1(n337), .A2(n2388), .B1(n2390), .B2(n137), .ZN(n1141) );
  OAI22_X2 U804 ( .A1(n336), .A2(n2388), .B1(n2390), .B2(n136), .ZN(n1140) );
  OAI22_X2 U805 ( .A1(n335), .A2(n2388), .B1(n2390), .B2(n135), .ZN(n1139) );
  OAI22_X2 U806 ( .A1(n380), .A2(n2388), .B1(n2390), .B2(n134), .ZN(n1138) );
  OAI22_X2 U807 ( .A1(n381), .A2(n2388), .B1(n2390), .B2(n133), .ZN(n1137) );
  OAI22_X2 U808 ( .A1(n379), .A2(n2388), .B1(n2390), .B2(n132), .ZN(n1136) );
  OAI22_X2 U809 ( .A1(n378), .A2(n2388), .B1(n2390), .B2(n131), .ZN(n1135) );
  OAI22_X2 U810 ( .A1(n377), .A2(n2388), .B1(n2390), .B2(n130), .ZN(n1134) );
  OAI22_X2 U811 ( .A1(n376), .A2(n2388), .B1(n2391), .B2(n129), .ZN(n1133) );
  OAI22_X2 U812 ( .A1(n375), .A2(n2389), .B1(n2391), .B2(n128), .ZN(n1132) );
  OAI22_X2 U813 ( .A1(n374), .A2(n2389), .B1(n2391), .B2(n127), .ZN(n1131) );
  OAI22_X2 U814 ( .A1(n373), .A2(n2389), .B1(n2391), .B2(n126), .ZN(n1130) );
  OAI22_X2 U815 ( .A1(n372), .A2(n2389), .B1(n2391), .B2(n125), .ZN(n1129) );
  OAI22_X2 U816 ( .A1(n370), .A2(n2389), .B1(n2391), .B2(n124), .ZN(n1128) );
  OAI22_X2 U817 ( .A1(n535), .A2(n2389), .B1(n2391), .B2(n123), .ZN(n1127) );
  OAI22_X2 U818 ( .A1(n384), .A2(n2389), .B1(n2391), .B2(n122), .ZN(n1126) );
  OAI22_X2 U819 ( .A1(n534), .A2(n2389), .B1(n2391), .B2(n121), .ZN(n1125) );
  OAI22_X2 U820 ( .A1(n2334), .A2(n2389), .B1(n2390), .B2(n119), .ZN(n1124) );
  NAND2_X2 U821 ( .A1(n610), .A2(n2387), .ZN(n966) );
  NAND4_X2 U824 ( .A1(n2022), .A2(n1590), .A3(n241), .A4(n240), .ZN(n915) );
  OAI22_X2 U825 ( .A1(n43), .A2(n69), .B1(n109), .B2(n1591), .ZN(n1113) );
  NAND2_X2 U826 ( .A1(n2435), .A2(n754), .ZN(n1591) );
  OAI22_X2 U827 ( .A1(n949), .A2(n1592), .B1(n900), .B2(n1593), .ZN(n1111) );
  XOR2_X2 U828 ( .A(n395), .B(n1594), .Z(n900) );
  OAI22_X2 U829 ( .A1(n948), .A2(n1592), .B1(n280), .B2(n1593), .ZN(n1110) );
  XOR2_X2 U830 ( .A(n282), .B(n1500), .Z(n1123) );
  OAI22_X2 U831 ( .A1(n947), .A2(n1592), .B1(n278), .B2(n1593), .ZN(n1109) );
  XNOR2_X2 U832 ( .A(n1595), .B(n1502), .ZN(n1299) );
  NAND2_X2 U833 ( .A1(n1596), .A2(n1597), .ZN(n1595) );
  OAI22_X2 U834 ( .A1(n946), .A2(n1592), .B1(n902), .B2(n1593), .ZN(n1108) );
  XOR2_X2 U835 ( .A(n277), .B(n1598), .Z(n902) );
  OAI22_X2 U836 ( .A1(n945), .A2(n1592), .B1(n903), .B2(n1593), .ZN(n1107) );
  XOR2_X2 U837 ( .A(n1600), .B(n1601), .Z(n903) );
  OAI22_X2 U840 ( .A1(n944), .A2(n1592), .B1(n271), .B2(n1593), .ZN(n1106) );
  NAND2_X2 U841 ( .A1(n41), .A2(n1592), .ZN(n1593) );
  XOR2_X2 U842 ( .A(n1315), .B(n1316), .Z(n1310) );
  XNOR2_X2 U843 ( .A(reg_a[5]), .B(reg_b[5]), .ZN(n1316) );
  OAI22_X2 U846 ( .A1(n274), .A2(n491), .B1(n1601), .B2(n1602), .ZN(n1539) );
  NAND2_X2 U847 ( .A1(reg_b[3]), .A2(reg_a[3]), .ZN(n1602) );
  OAI22_X2 U848 ( .A1(n279), .A2(n492), .B1(n1502), .B2(n1596), .ZN(n1603) );
  NAND2_X2 U849 ( .A1(reg_b[1]), .A2(reg_a[1]), .ZN(n1596) );
  XOR2_X2 U851 ( .A(reg_a[2]), .B(n279), .Z(n1502) );
  NAND2_X2 U852 ( .A1(n1500), .A2(n282), .ZN(n1597) );
  AOI22_X2 U853 ( .A1(n1594), .A2(reg_carry), .B1(reg_a[0]), .B2(reg_b[0]), 
        .ZN(n1501) );
  XOR2_X2 U854 ( .A(reg_a[0]), .B(reg_b[0]), .Z(n1594) );
  XOR2_X2 U855 ( .A(reg_a[1]), .B(reg_b[1]), .Z(n1500) );
  XOR2_X2 U857 ( .A(n491), .B(reg_b[4]), .Z(n1601) );
  XNOR2_X2 U858 ( .A(reg_a[3]), .B(reg_b[3]), .ZN(n1598) );
  NAND2_X2 U860 ( .A1(n107), .A2(n968), .ZN(n901) );
  OAI22_X2 U861 ( .A1(n3285), .A2(n1605), .B1(n100), .B2(n2369), .ZN(n1105) );
  OAI22_X2 U862 ( .A1(n3284), .A2(n1607), .B1(n99), .B2(n2369), .ZN(n1104) );
  OAI22_X2 U863 ( .A1(n1608), .A2(n218), .B1(n98), .B2(n2369), .ZN(n1103) );
  OAI22_X2 U864 ( .A1(n1609), .A2(n216), .B1(n97), .B2(n2369), .ZN(n1102) );
  OAI22_X2 U865 ( .A1(n1610), .A2(n215), .B1(n96), .B2(n2369), .ZN(n1101) );
  OAI22_X2 U866 ( .A1(n1611), .A2(n214), .B1(n95), .B2(n2369), .ZN(n1100) );
  OAI22_X2 U867 ( .A1(n1612), .A2(n213), .B1(n94), .B2(n2369), .ZN(n1099) );
  OAI22_X2 U868 ( .A1(n1613), .A2(n219), .B1(n93), .B2(n2369), .ZN(n1098) );
  OAI22_X2 U869 ( .A1(n1614), .A2(n235), .B1(n92), .B2(n2369), .ZN(n1097) );
  OAI22_X2 U870 ( .A1(n1615), .A2(n234), .B1(n91), .B2(n2368), .ZN(n1096) );
  OAI22_X2 U871 ( .A1(n1616), .A2(n233), .B1(n90), .B2(n2368), .ZN(n1095) );
  OAI22_X2 U872 ( .A1(n1617), .A2(n232), .B1(n89), .B2(n2368), .ZN(n1094) );
  OAI22_X2 U873 ( .A1(n1618), .A2(n231), .B1(n88), .B2(n2368), .ZN(n1093) );
  OAI22_X2 U874 ( .A1(n1619), .A2(n230), .B1(n87), .B2(n2368), .ZN(n1092) );
  OAI22_X2 U875 ( .A1(n1620), .A2(n229), .B1(n86), .B2(n2368), .ZN(n1091) );
  OAI22_X2 U876 ( .A1(n1621), .A2(n228), .B1(n85), .B2(n2368), .ZN(n1090) );
  OAI22_X2 U877 ( .A1(n1622), .A2(n227), .B1(n84), .B2(n2368), .ZN(n1089) );
  OAI22_X2 U878 ( .A1(n1623), .A2(n226), .B1(n83), .B2(n2368), .ZN(n1088) );
  OAI22_X2 U879 ( .A1(n1624), .A2(n225), .B1(n82), .B2(n2368), .ZN(n1087) );
  OAI22_X2 U880 ( .A1(n1625), .A2(n224), .B1(n81), .B2(n2368), .ZN(n1086) );
  OAI22_X2 U881 ( .A1(n1626), .A2(n223), .B1(n80), .B2(n2367), .ZN(n1085) );
  OAI22_X2 U882 ( .A1(n1627), .A2(n222), .B1(n79), .B2(n2367), .ZN(n1084) );
  OAI22_X2 U883 ( .A1(n1628), .A2(n221), .B1(n78), .B2(n2367), .ZN(n1083) );
  OAI22_X2 U884 ( .A1(n1629), .A2(n220), .B1(n77), .B2(n2367), .ZN(n1082) );
  OAI22_X2 U885 ( .A1(n1630), .A2(n189), .B1(n76), .B2(n2367), .ZN(n1081) );
  OAI22_X2 U886 ( .A1(n1631), .A2(n188), .B1(n75), .B2(n2367), .ZN(n1080) );
  OAI22_X2 U887 ( .A1(n1632), .A2(n187), .B1(n74), .B2(n2367), .ZN(n1079) );
  OAI22_X2 U888 ( .A1(n1633), .A2(n186), .B1(n73), .B2(n2367), .ZN(n1078) );
  OAI22_X2 U889 ( .A1(n1634), .A2(n185), .B1(n72), .B2(n2367), .ZN(n1077) );
  OAI22_X2 U890 ( .A1(n1635), .A2(n184), .B1(n71), .B2(n2367), .ZN(n1076) );
  OAI22_X2 U891 ( .A1(n1636), .A2(n183), .B1(n70), .B2(n2367), .ZN(n1075) );
  OAI22_X2 U893 ( .A1(n100), .A2(n2366), .B1(n398), .B2(n1605), .ZN(n1074) );
  OAI22_X2 U895 ( .A1(n99), .A2(n2366), .B1(n195), .B2(n1607), .ZN(n1073) );
  OAI22_X2 U897 ( .A1(n98), .A2(n2366), .B1(n194), .B2(n1608), .ZN(n1072) );
  OAI22_X2 U899 ( .A1(n97), .A2(n2366), .B1(n193), .B2(n1609), .ZN(n1071) );
  OAI22_X2 U901 ( .A1(n96), .A2(n2366), .B1(n192), .B2(n1610), .ZN(n1070) );
  OAI22_X2 U903 ( .A1(n95), .A2(n2366), .B1(n196), .B2(n1611), .ZN(n1069) );
  OAI22_X2 U905 ( .A1(n94), .A2(n2366), .B1(n191), .B2(n1612), .ZN(n1068) );
  OAI22_X2 U907 ( .A1(n93), .A2(n2366), .B1(n190), .B2(n1613), .ZN(n1067) );
  OAI22_X2 U910 ( .A1(n92), .A2(n2366), .B1(n200), .B2(n1614), .ZN(n1066) );
  OAI22_X2 U912 ( .A1(n91), .A2(n2365), .B1(n199), .B2(n1615), .ZN(n1065) );
  OAI22_X2 U914 ( .A1(n90), .A2(n2365), .B1(n198), .B2(n1616), .ZN(n1064) );
  OAI22_X2 U916 ( .A1(n89), .A2(n2365), .B1(n197), .B2(n1617), .ZN(n1063) );
  OAI22_X2 U918 ( .A1(n88), .A2(n2365), .B1(n212), .B2(n1618), .ZN(n1062) );
  OAI22_X2 U920 ( .A1(n87), .A2(n2365), .B1(n211), .B2(n1619), .ZN(n1061) );
  OAI22_X2 U922 ( .A1(n86), .A2(n2365), .B1(n210), .B2(n1620), .ZN(n1060) );
  OAI22_X2 U924 ( .A1(n85), .A2(n2365), .B1(n209), .B2(n1621), .ZN(n1059) );
  OAI22_X2 U927 ( .A1(n84), .A2(n2365), .B1(n208), .B2(n1622), .ZN(n1058) );
  OAI22_X2 U929 ( .A1(n83), .A2(n2365), .B1(n207), .B2(n1623), .ZN(n1057) );
  OAI22_X2 U931 ( .A1(n82), .A2(n2365), .B1(n206), .B2(n1624), .ZN(n1056) );
  OAI22_X2 U933 ( .A1(n81), .A2(n2365), .B1(n205), .B2(n1625), .ZN(n1055) );
  OAI22_X2 U935 ( .A1(n80), .A2(n2364), .B1(n204), .B2(n1626), .ZN(n1054) );
  OAI22_X2 U937 ( .A1(n79), .A2(n2364), .B1(n203), .B2(n1627), .ZN(n1053) );
  OAI22_X2 U939 ( .A1(n78), .A2(n2364), .B1(n202), .B2(n1628), .ZN(n1052) );
  OAI22_X2 U941 ( .A1(n77), .A2(n2364), .B1(n201), .B2(n1629), .ZN(n1051) );
  OAI22_X2 U945 ( .A1(n76), .A2(n2364), .B1(n181), .B2(n1630), .ZN(n1050) );
  OAI22_X2 U948 ( .A1(n75), .A2(n2364), .B1(n180), .B2(n1631), .ZN(n1049) );
  OAI22_X2 U951 ( .A1(n74), .A2(n2364), .B1(n179), .B2(n1632), .ZN(n1048) );
  OAI22_X2 U954 ( .A1(n73), .A2(n2364), .B1(n178), .B2(n1633), .ZN(n1047) );
  OAI22_X2 U957 ( .A1(n72), .A2(n2364), .B1(n177), .B2(n1634), .ZN(n1046) );
  OAI22_X2 U960 ( .A1(n71), .A2(n2364), .B1(n176), .B2(n1635), .ZN(n1045) );
  OAI22_X2 U963 ( .A1(n182), .A2(n1636), .B1(n70), .B2(n2364), .ZN(n1044) );
  NAND4_X2 U967 ( .A1(state[0]), .A2(n1651), .A3(n239), .A4(n238), .ZN(n913)
         );
  NAND4_X2 U970 ( .A1(state[2]), .A2(n1651), .A3(n105), .A4(n239), .ZN(n611)
         );
  OAI211_X2 U972 ( .C1(n2419), .C2(n395), .A(n1652), .B(n899), .ZN(n1043) );
  NAND4_X2 U975 ( .A1(n1654), .A2(n1655), .A3(n1656), .A4(n1657), .ZN(n1042)
         );
  AOI22_X2 U976 ( .A1(n40), .A2(n1950), .B1(n2360), .B2(n399), .ZN(n1657) );
  AOI22_X2 U977 ( .A1(n3285), .A2(n2026), .B1(n2359), .B2(i_divisor[0]), .ZN(
        n1656) );
  AOI22_X2 U978 ( .A1(n2354), .A2(n580), .B1(n2353), .B2(n118), .ZN(n1655) );
  AOI22_X2 U979 ( .A1(n2350), .A2(n3187), .B1(reg_a[0]), .B2(n2416), .ZN(n1654) );
  NAND4_X2 U980 ( .A1(n1664), .A2(n1665), .A3(n1666), .A4(n1667), .ZN(n1041)
         );
  AOI22_X2 U983 ( .A1(n40), .A2(n1953), .B1(n2359), .B2(i_divisor[1]), .ZN(
        n1666) );
  AOI22_X2 U984 ( .A1(n2354), .A2(n579), .B1(n2353), .B2(n117), .ZN(n1665) );
  AOI22_X2 U985 ( .A1(n2350), .A2(n3122), .B1(reg_a[1]), .B2(n2417), .ZN(n1664) );
  NAND4_X2 U986 ( .A1(n1670), .A2(n1671), .A3(n1672), .A4(n1673), .ZN(n1040)
         );
  AOI22_X2 U987 ( .A1(n20), .A2(n218), .B1(n40), .B2(n1952), .ZN(n1673) );
  AOI22_X2 U990 ( .A1(n1675), .A2(n2362), .B1(n2359), .B2(i_divisor[2]), .ZN(
        n1672) );
  AOI22_X2 U991 ( .A1(n2354), .A2(n578), .B1(n2353), .B2(n116), .ZN(n1671) );
  AOI22_X2 U992 ( .A1(n2350), .A2(n3125), .B1(reg_a[2]), .B2(n2416), .ZN(n1670) );
  NAND4_X2 U993 ( .A1(n1676), .A2(n1677), .A3(n1678), .A4(n1679), .ZN(n1039)
         );
  AOI22_X2 U996 ( .A1(n40), .A2(n1951), .B1(n2359), .B2(i_divisor[3]), .ZN(
        n1678) );
  NAND2_X2 U997 ( .A1(n1976), .A2(n2419), .ZN(n756) );
  AOI22_X2 U998 ( .A1(n2354), .A2(n577), .B1(n2353), .B2(n115), .ZN(n1677) );
  AOI22_X2 U999 ( .A1(n2350), .A2(n3128), .B1(reg_a[3]), .B2(n2416), .ZN(n1676) );
  AOI22_X2 U1002 ( .A1(n19), .A2(n215), .B1(n1685), .B2(n2362), .ZN(n1683) );
  AOI22_X2 U1005 ( .A1(n2359), .A2(i_divisor[4]), .B1(n2354), .B2(n576), .ZN(
        n1682) );
  NAND4_X2 U1006 ( .A1(n1687), .A2(n1688), .A3(n1689), .A4(n1690), .ZN(n1037)
         );
  AOI22_X2 U1008 ( .A1(n2359), .A2(i_divisor[5]), .B1(n2356), .B2(n575), .ZN(
        n1689) );
  NAND2_X2 U1010 ( .A1(n1691), .A2(n214), .ZN(n1687) );
  AOI22_X2 U1013 ( .A1(n1695), .A2(n213), .B1(n1696), .B2(n2362), .ZN(n1693)
         );
  AOI22_X2 U1016 ( .A1(n2359), .A2(i_divisor[6]), .B1(n2356), .B2(n574), .ZN(
        n1692) );
  NAND4_X2 U1017 ( .A1(n1697), .A2(n1698), .A3(n1699), .A4(n1700), .ZN(n1035)
         );
  AOI22_X2 U1019 ( .A1(n2359), .A2(i_divisor[7]), .B1(n2356), .B2(n573), .ZN(
        n1699) );
  NAND2_X2 U1021 ( .A1(n1701), .A2(n219), .ZN(n1697) );
  AOI22_X2 U1024 ( .A1(n1705), .A2(n235), .B1(n1706), .B2(n2362), .ZN(n1703)
         );
  AOI22_X2 U1027 ( .A1(n2358), .A2(i_divisor[8]), .B1(n2356), .B2(n572), .ZN(
        n1702) );
  NAND4_X2 U1028 ( .A1(n1707), .A2(n1708), .A3(n1709), .A4(n1710), .ZN(n1033)
         );
  AOI22_X2 U1030 ( .A1(n2358), .A2(i_divisor[9]), .B1(n2356), .B2(n571), .ZN(
        n1709) );
  NAND2_X2 U1032 ( .A1(n1711), .A2(n234), .ZN(n1707) );
  AOI22_X2 U1035 ( .A1(n1715), .A2(n233), .B1(n1716), .B2(n2362), .ZN(n1713)
         );
  AOI22_X2 U1038 ( .A1(n2358), .A2(i_divisor[10]), .B1(n2356), .B2(n570), .ZN(
        n1712) );
  NAND4_X2 U1039 ( .A1(n1717), .A2(n1718), .A3(n1719), .A4(n1720), .ZN(n1031)
         );
  AOI22_X2 U1041 ( .A1(n2358), .A2(i_divisor[11]), .B1(n2356), .B2(n569), .ZN(
        n1719) );
  NAND2_X2 U1043 ( .A1(n1721), .A2(n232), .ZN(n1717) );
  AOI22_X2 U1046 ( .A1(n1725), .A2(n231), .B1(n1726), .B2(n2362), .ZN(n1723)
         );
  AOI22_X2 U1049 ( .A1(n2358), .A2(i_divisor[12]), .B1(n2356), .B2(n568), .ZN(
        n1722) );
  NAND4_X2 U1050 ( .A1(n1727), .A2(n1728), .A3(n1729), .A4(n1730), .ZN(n1029)
         );
  AOI22_X2 U1052 ( .A1(n2358), .A2(i_divisor[13]), .B1(n2355), .B2(n567), .ZN(
        n1729) );
  NAND2_X2 U1054 ( .A1(n1731), .A2(n230), .ZN(n1727) );
  AOI22_X2 U1057 ( .A1(n1735), .A2(n229), .B1(n1736), .B2(n2362), .ZN(n1733)
         );
  AOI22_X2 U1060 ( .A1(n2358), .A2(i_divisor[14]), .B1(n2355), .B2(n566), .ZN(
        n1732) );
  NAND4_X2 U1061 ( .A1(n1737), .A2(n1738), .A3(n1739), .A4(n1740), .ZN(n1027)
         );
  AOI22_X2 U1063 ( .A1(n2358), .A2(i_divisor[15]), .B1(n2355), .B2(n565), .ZN(
        n1739) );
  NAND2_X2 U1065 ( .A1(n1741), .A2(n228), .ZN(n1737) );
  AOI22_X2 U1068 ( .A1(n1745), .A2(n227), .B1(n1746), .B2(n2362), .ZN(n1743)
         );
  AOI22_X2 U1071 ( .A1(n2358), .A2(i_divisor[16]), .B1(n2355), .B2(n564), .ZN(
        n1742) );
  NAND4_X2 U1072 ( .A1(n1747), .A2(n1748), .A3(n1749), .A4(n1750), .ZN(n1025)
         );
  AOI22_X2 U1074 ( .A1(n2358), .A2(i_divisor[17]), .B1(n2355), .B2(n563), .ZN(
        n1749) );
  NAND2_X2 U1076 ( .A1(n1751), .A2(n226), .ZN(n1747) );
  AOI22_X2 U1079 ( .A1(n1755), .A2(n225), .B1(n1756), .B2(n2362), .ZN(n1753)
         );
  AOI22_X2 U1082 ( .A1(n2358), .A2(i_divisor[18]), .B1(n2355), .B2(n562), .ZN(
        n1752) );
  NAND4_X2 U1083 ( .A1(n1757), .A2(n1758), .A3(n1759), .A4(n1760), .ZN(n1023)
         );
  AOI22_X2 U1085 ( .A1(n2358), .A2(i_divisor[19]), .B1(n2355), .B2(n561), .ZN(
        n1759) );
  NAND2_X2 U1087 ( .A1(n1761), .A2(n224), .ZN(n1757) );
  AOI22_X2 U1090 ( .A1(n1765), .A2(n223), .B1(n1766), .B2(n2362), .ZN(n1763)
         );
  AOI22_X2 U1093 ( .A1(n2357), .A2(i_divisor[20]), .B1(n2355), .B2(n560), .ZN(
        n1762) );
  NAND4_X2 U1094 ( .A1(n1767), .A2(n1768), .A3(n1769), .A4(n1770), .ZN(n1021)
         );
  AOI22_X2 U1096 ( .A1(n2357), .A2(i_divisor[21]), .B1(n2355), .B2(n559), .ZN(
        n1769) );
  NAND2_X2 U1098 ( .A1(n1771), .A2(n222), .ZN(n1767) );
  AOI22_X2 U1101 ( .A1(n1775), .A2(n221), .B1(n1776), .B2(n2362), .ZN(n1773)
         );
  AOI22_X2 U1104 ( .A1(n2357), .A2(i_divisor[22]), .B1(n2355), .B2(n558), .ZN(
        n1772) );
  NAND4_X2 U1105 ( .A1(n1777), .A2(n1778), .A3(n1779), .A4(n1780), .ZN(n1019)
         );
  AOI22_X2 U1107 ( .A1(n2357), .A2(i_divisor[23]), .B1(n2355), .B2(n557), .ZN(
        n1779) );
  NAND2_X2 U1109 ( .A1(n1781), .A2(n220), .ZN(n1777) );
  AOI22_X2 U1112 ( .A1(n1785), .A2(n2362), .B1(n9), .B2(n189), .ZN(n1783) );
  AOI22_X2 U1113 ( .A1(n2357), .A2(i_divisor[24]), .B1(n2355), .B2(n556), .ZN(
        n1782) );
  AOI22_X2 U1116 ( .A1(n1790), .A2(n188), .B1(n1791), .B2(n2362), .ZN(n1788)
         );
  AOI22_X2 U1120 ( .A1(n2357), .A2(i_divisor[25]), .B1(n2354), .B2(n555), .ZN(
        n1787) );
  NAND4_X2 U1121 ( .A1(n1792), .A2(n1793), .A3(n1794), .A4(n1795), .ZN(n1016)
         );
  AOI22_X2 U1123 ( .A1(n2357), .A2(i_divisor[26]), .B1(n2354), .B2(n554), .ZN(
        n1794) );
  NAND2_X2 U1125 ( .A1(n1796), .A2(n187), .ZN(n1792) );
  AOI22_X2 U1128 ( .A1(n1800), .A2(n2362), .B1(n8), .B2(n186), .ZN(n1798) );
  AOI22_X2 U1129 ( .A1(n2357), .A2(i_divisor[27]), .B1(n2354), .B2(n553), .ZN(
        n1797) );
  AOI22_X2 U1132 ( .A1(n1805), .A2(n185), .B1(n1806), .B2(n2362), .ZN(n1803)
         );
  AOI22_X2 U1136 ( .A1(n2357), .A2(i_divisor[28]), .B1(n2354), .B2(n552), .ZN(
        n1802) );
  NAND4_X2 U1137 ( .A1(n1807), .A2(n1808), .A3(n1809), .A4(n1810), .ZN(n1013)
         );
  AOI22_X2 U1139 ( .A1(n2357), .A2(i_divisor[29]), .B1(n2354), .B2(n551), .ZN(
        n1809) );
  NAND2_X2 U1140 ( .A1(n1811), .A2(n184), .ZN(n1807) );
  OAI22_X2 U1143 ( .A1(n1815), .A2(nq[30]), .B1(n1808), .B2(n183), .ZN(n1814)
         );
  AND2_X2 U1148 ( .A1(n1800), .A2(nq[28]), .ZN(n1806) );
  AND3_X2 U1149 ( .A1(nq[27]), .A2(nq[26]), .A3(n1791), .ZN(n1800) );
  AND2_X2 U1150 ( .A1(n1785), .A2(nq[25]), .ZN(n1791) );
  AND3_X2 U1151 ( .A1(nq[24]), .A2(nq[23]), .A3(n1776), .ZN(n1785) );
  AND3_X2 U1152 ( .A1(nq[22]), .A2(nq[21]), .A3(n1766), .ZN(n1776) );
  AND3_X2 U1153 ( .A1(nq[20]), .A2(nq[19]), .A3(n1756), .ZN(n1766) );
  AND3_X2 U1154 ( .A1(nq[18]), .A2(nq[17]), .A3(n1746), .ZN(n1756) );
  AND3_X2 U1155 ( .A1(nq[16]), .A2(nq[15]), .A3(n1736), .ZN(n1746) );
  AND3_X2 U1156 ( .A1(nq[14]), .A2(nq[13]), .A3(n1726), .ZN(n1736) );
  AND3_X2 U1157 ( .A1(nq[12]), .A2(nq[11]), .A3(n1716), .ZN(n1726) );
  AND3_X2 U1158 ( .A1(nq[10]), .A2(nq[9]), .A3(n1706), .ZN(n1716) );
  AND3_X2 U1159 ( .A1(nq[8]), .A2(nq[7]), .A3(n1696), .ZN(n1706) );
  AND3_X2 U1160 ( .A1(nq[6]), .A2(nq[5]), .A3(n1685), .ZN(n1696) );
  AOI22_X2 U1164 ( .A1(n2357), .A2(i_divisor[30]), .B1(n2354), .B2(n550), .ZN(
        n1812) );
  NAND2_X2 U1165 ( .A1(n1817), .A2(n1818), .ZN(n1011) );
  AOI221_X2 U1166 ( .B1(n2354), .B2(n549), .C1(n2357), .C2(i_divisor[31]), .A(
        n37), .ZN(n1818) );
  XOR2_X2 U1173 ( .A(n1955), .B(n284), .Z(n1819) );
  NAND2_X2 U1174 ( .A1(n1821), .A2(n1822), .ZN(n1820) );
  NOR4_X2 U1175 ( .A1(n1823), .A2(n1824), .A3(n1825), .A4(n1826), .ZN(n1822)
         );
  NAND4_X2 U1176 ( .A1(n151), .A2(n156), .A3(n168), .A4(n155), .ZN(n1826) );
  NAND4_X2 U1177 ( .A1(n165), .A2(n164), .A3(n166), .A4(n167), .ZN(n1825) );
  NAND4_X2 U1178 ( .A1(n153), .A2(n152), .A3(n158), .A4(n157), .ZN(n1824) );
  NAND4_X2 U1179 ( .A1(n163), .A2(n161), .A3(n160), .A4(n159), .ZN(n1823) );
  NOR4_X2 U1180 ( .A1(n1827), .A2(n1828), .A3(n1829), .A4(n1830), .ZN(n1821)
         );
  OR4_X2 U1181 ( .A1(n284), .A2(n3053), .A3(n3120), .A4(n3123), .ZN(n1830) );
  OR4_X2 U1182 ( .A1(n3126), .A2(n3129), .A3(n3132), .A4(n1977), .ZN(n1829) );
  NAND4_X2 U1183 ( .A1(n149), .A2(n144), .A3(n148), .A4(n162), .ZN(n1828) );
  NAND4_X2 U1184 ( .A1(n150), .A2(n147), .A3(n146), .A4(n145), .ZN(n1827) );
  XNOR2_X2 U1188 ( .A(n284), .B(n3193), .ZN(n1650) );
  NAND4_X2 U1189 ( .A1(n964), .A2(n963), .A3(n2418), .A4(n109), .ZN(n757) );
  NAND4_X2 U1190 ( .A1(state[4]), .A2(n1590), .A3(n241), .A4(n2335), .ZN(n964)
         );
  NAND2_X2 U1192 ( .A1(state_reg_1_0), .A2(n110), .ZN(n612) );
  NAND2_X2 U1193 ( .A1(n1831), .A2(n1832), .ZN(n1010) );
  AOI221_X2 U1194 ( .B1(n2339), .B2(n1833), .C1(n641), .C2(n1834), .A(n1835), 
        .ZN(n1832) );
  OAI221_X2 U1195 ( .B1(n411), .B2(n666), .C1(n430), .C2(n63), .A(n668), .ZN(
        n1835) );
  OAI221_X2 U1196 ( .B1(n429), .B2(n672), .C1(n426), .C2(n1836), .A(n1837), 
        .ZN(n682) );
  AOI22_X2 U1197 ( .A1(n1838), .A2(n650), .B1(n1839), .B2(n651), .ZN(n1837) );
  AOI221_X2 U1198 ( .B1(n2430), .B2(sdata[0]), .C1(i_dividend[0]), .C2(n2426), 
        .A(n1840), .ZN(n1831) );
  OAI22_X2 U1199 ( .A1(n1978), .A2(n2337), .B1(n1841), .B2(n2024), .ZN(n1840)
         );
  AOI221_X2 U1200 ( .B1(n2016), .B2(n466), .C1(n2018), .C2(n478), .A(n1842), 
        .ZN(n1841) );
  OAI22_X2 U1201 ( .A1(n1984), .A2(n1843), .B1(n1980), .B2(n1844), .ZN(n1842)
         );
  OAI221_X2 U1202 ( .B1(n1845), .B2(n719), .C1(n1979), .C2(n2337), .A(n1846), 
        .ZN(n1009) );
  AOI22_X2 U1203 ( .A1(n2431), .A2(sdata[1]), .B1(i_dividend[1]), .B2(n2427), 
        .ZN(n1846) );
  OAI22_X2 U1205 ( .A1(n424), .A2(n1850), .B1(n1851), .B2(n405), .ZN(n1849) );
  OAI221_X2 U1206 ( .B1(n1852), .B2(n1853), .C1(n1854), .C2(n1855), .A(n1856), 
        .ZN(n1848) );
  AOI221_X2 U1207 ( .B1(n2016), .B2(n478), .C1(n2018), .C2(n473), .A(n1857), 
        .ZN(n1854) );
  OAI22_X2 U1208 ( .A1(n1980), .A2(n1843), .B1(n1985), .B2(n1844), .ZN(n1857)
         );
  AOI221_X2 U1209 ( .B1(n1838), .B2(n440), .C1(n1839), .C2(n659), .A(n1858), 
        .ZN(n1852) );
  OAI22_X2 U1210 ( .A1(n421), .A2(n1836), .B1(n423), .B2(n672), .ZN(n1858) );
  OAI221_X2 U1211 ( .B1(n1859), .B2(n719), .C1(n1984), .C2(n2336), .A(n1860), 
        .ZN(n1008) );
  AOI22_X2 U1212 ( .A1(n2430), .A2(sdata[2]), .B1(i_dividend[2]), .B2(n2427), 
        .ZN(n1860) );
  OAI22_X2 U1214 ( .A1(n419), .A2(n1850), .B1(n1865), .B2(n405), .ZN(n1863) );
  OAI221_X2 U1215 ( .B1(n1866), .B2(n1853), .C1(n1867), .C2(n1855), .A(n1856), 
        .ZN(n1862) );
  AOI221_X2 U1216 ( .B1(n2016), .B2(n473), .C1(n2018), .C2(n477), .A(n1868), 
        .ZN(n1867) );
  OAI22_X2 U1217 ( .A1(n1985), .A2(n1843), .B1(n1986), .B2(n1844), .ZN(n1868)
         );
  AOI221_X2 U1218 ( .B1(n1838), .B2(n670), .C1(n1839), .C2(n671), .A(n690), 
        .ZN(n1866) );
  OAI22_X2 U1219 ( .A1(n418), .A2(n672), .B1(n416), .B2(n1836), .ZN(n690) );
  OAI221_X2 U1220 ( .B1(n1870), .B2(n719), .C1(n1980), .C2(n634), .A(n1871), 
        .ZN(n1007) );
  AOI22_X2 U1221 ( .A1(sdata[3]), .A2(n2431), .B1(i_dividend[3]), .B2(n2427), 
        .ZN(n1871) );
  OAI22_X2 U1223 ( .A1(n435), .A2(n1850), .B1(n436), .B2(n1869), .ZN(n1875) );
  OAI221_X2 U1224 ( .B1(n410), .B2(n1853), .C1(n1876), .C2(n1855), .A(n1856), 
        .ZN(n1874) );
  AOI221_X2 U1225 ( .B1(n2016), .B2(n477), .C1(n2018), .C2(n472), .A(n1877), 
        .ZN(n1876) );
  OAI22_X2 U1226 ( .A1(n1986), .A2(n1843), .B1(n1987), .B2(n1844), .ZN(n1877)
         );
  OAI221_X2 U1227 ( .B1(n1836), .B2(n433), .C1(n672), .C2(n432), .A(n1879), 
        .ZN(n1878) );
  NAND2_X2 U1229 ( .A1(n1880), .A2(n1881), .ZN(n1006) );
  AOI221_X2 U1230 ( .B1(n2339), .B2(n653), .C1(n641), .C2(n1833), .A(n1882), 
        .ZN(n1881) );
  OAI221_X2 U1231 ( .B1(n409), .B2(n666), .C1(n429), .C2(n63), .A(n668), .ZN(
        n1882) );
  OAI221_X2 U1232 ( .B1(n427), .B2(n1836), .C1(n426), .C2(n672), .A(n1883), 
        .ZN(n698) );
  AOI221_X2 U1234 ( .B1(sdata[4]), .B2(n2430), .C1(i_dividend[4]), .C2(n2426), 
        .A(n1884), .ZN(n1880) );
  OAI22_X2 U1235 ( .A1(n1985), .A2(n2336), .B1(n437), .B2(n2024), .ZN(n1884)
         );
  OAI221_X2 U1236 ( .B1(n1985), .B2(n2347), .C1(n1986), .C2(n2345), .A(n1887), 
        .ZN(n1834) );
  AOI22_X2 U1237 ( .A1(n438), .A2(n469), .B1(n439), .B2(n470), .ZN(n1887) );
  NAND2_X2 U1238 ( .A1(n1888), .A2(n1889), .ZN(n1005) );
  AOI221_X2 U1239 ( .B1(n2339), .B2(n661), .C1(n641), .C2(n1847), .A(n1890), 
        .ZN(n1889) );
  OAI221_X2 U1240 ( .B1(n408), .B2(n666), .C1(n423), .C2(n63), .A(n668), .ZN(
        n1890) );
  OAI221_X2 U1241 ( .B1(n422), .B2(n1836), .C1(n421), .C2(n672), .A(n1891), 
        .ZN(n700) );
  AOI221_X2 U1243 ( .B1(sdata[5]), .B2(n2430), .C1(i_dividend[5]), .C2(n2426), 
        .A(n1892), .ZN(n1888) );
  OAI22_X2 U1244 ( .A1(n1986), .A2(n2337), .B1(n1851), .B2(n2024), .ZN(n1892)
         );
  AOI221_X2 U1245 ( .B1(n471), .B2(n2016), .C1(n470), .C2(n2018), .A(n1893), 
        .ZN(n1851) );
  OAI22_X2 U1246 ( .A1(n1844), .A2(n1989), .B1(n1843), .B2(n1988), .ZN(n1893)
         );
  NAND2_X2 U1247 ( .A1(n1894), .A2(n1895), .ZN(n1004) );
  AOI221_X2 U1248 ( .B1(n2339), .B2(n674), .C1(n641), .C2(n1861), .A(n1896), 
        .ZN(n1895) );
  OAI221_X2 U1249 ( .B1(n407), .B2(n666), .C1(n418), .C2(n63), .A(n668), .ZN(
        n1896) );
  NAND2_X2 U1250 ( .A1(n400), .A2(n2425), .ZN(n668) );
  NAND2_X2 U1252 ( .A1(n402), .A2(n2425), .ZN(n666) );
  OAI221_X2 U1253 ( .B1(n417), .B2(n1836), .C1(n416), .C2(n672), .A(n1897), 
        .ZN(n702) );
  AND2_X2 U1255 ( .A1(n712), .A2(n414), .ZN(n694) );
  AOI221_X2 U1258 ( .B1(sdata[6]), .B2(n2430), .C1(i_dividend[6]), .C2(n2426), 
        .A(n1898), .ZN(n1894) );
  OAI22_X2 U1259 ( .A1(n1987), .A2(n2336), .B1(n1865), .B2(n2024), .ZN(n1898)
         );
  AOI221_X2 U1261 ( .B1(n470), .B2(n2016), .C1(n469), .C2(n2018), .A(n1899), 
        .ZN(n1865) );
  OAI22_X2 U1262 ( .A1(n1844), .A2(n1990), .B1(n1843), .B2(n1989), .ZN(n1899)
         );
  OAI221_X2 U1263 ( .B1(n1900), .B2(n719), .C1(n1988), .C2(n2337), .A(n1901), 
        .ZN(n1003) );
  AOI22_X2 U1264 ( .A1(sdata[7]), .A2(n2431), .B1(i_dividend[7]), .B2(n2427), 
        .ZN(n1901) );
  OAI22_X2 U1266 ( .A1(n435), .A2(n1869), .B1(n436), .B2(n405), .ZN(n1904) );
  OAI221_X2 U1267 ( .B1(n2004), .B2(n2346), .C1(n2001), .C2(n2345), .A(n1905), 
        .ZN(n644) );
  AOI22_X2 U1268 ( .A1(n438), .A2(n448), .B1(n439), .B2(n449), .ZN(n1905) );
  OAI221_X2 U1269 ( .B1(n2002), .B2(n2346), .C1(n2007), .C2(n2345), .A(n1906), 
        .ZN(n642) );
  AOI22_X2 U1270 ( .A1(n438), .A2(n446), .B1(n439), .B2(n451), .ZN(n1906) );
  OAI22_X2 U1271 ( .A1(n433), .A2(n1907), .B1(n434), .B2(n1908), .ZN(n1903) );
  OAI221_X2 U1272 ( .B1(n1997), .B2(n2346), .C1(n1998), .C2(n2345), .A(n1909), 
        .ZN(n638) );
  AOI22_X2 U1273 ( .A1(n438), .A2(n456), .B1(n439), .B2(n457), .ZN(n1909) );
  OAI221_X2 U1274 ( .B1(n1993), .B2(n2346), .C1(n1994), .C2(n2345), .A(n1910), 
        .ZN(n640) );
  AOI22_X2 U1275 ( .A1(n438), .A2(n460), .B1(n439), .B2(n461), .ZN(n1910) );
  OAI221_X2 U1276 ( .B1(n431), .B2(n1855), .C1(n432), .C2(n1850), .A(n1911), 
        .ZN(n1902) );
  OAI221_X2 U1277 ( .B1(n1982), .B2(n2346), .C1(n1983), .C2(n2345), .A(n1912), 
        .ZN(n636) );
  AOI22_X2 U1278 ( .A1(n438), .A2(n464), .B1(n439), .B2(n465), .ZN(n1912) );
  OAI221_X2 U1279 ( .B1(n1988), .B2(n2346), .C1(n1989), .C2(n2345), .A(n1913), 
        .ZN(n1873) );
  AOI22_X2 U1280 ( .A1(n438), .A2(n476), .B1(n439), .B2(n467), .ZN(n1913) );
  OAI221_X2 U1281 ( .B1(n1914), .B2(n719), .C1(n1989), .C2(n2336), .A(n1915), 
        .ZN(n1002) );
  AOI22_X2 U1282 ( .A1(sdata[8]), .A2(n2431), .B1(i_dividend[8]), .B2(n2427), 
        .ZN(n1915) );
  OAI22_X2 U1284 ( .A1(n429), .A2(n1869), .B1(n430), .B2(n405), .ZN(n1918) );
  OAI221_X2 U1285 ( .B1(n2001), .B2(n2346), .C1(n2005), .C2(n2345), .A(n1919), 
        .ZN(n653) );
  AOI22_X2 U1286 ( .A1(n438), .A2(n452), .B1(n439), .B2(n448), .ZN(n1919) );
  OAI221_X2 U1287 ( .B1(n2007), .B2(n2346), .C1(n2003), .C2(n2345), .A(n1920), 
        .ZN(n652) );
  AOI22_X2 U1288 ( .A1(n438), .A2(n475), .B1(n439), .B2(n446), .ZN(n1920) );
  OAI22_X2 U1289 ( .A1(n427), .A2(n1907), .B1(n428), .B2(n1908), .ZN(n1917) );
  OAI221_X2 U1290 ( .B1(n1998), .B2(n2346), .C1(n1999), .C2(n2345), .A(n1921), 
        .ZN(n650) );
  AOI22_X2 U1291 ( .A1(n438), .A2(n455), .B1(n439), .B2(n456), .ZN(n1921) );
  OAI221_X2 U1292 ( .B1(n1994), .B2(n2346), .C1(n1995), .C2(n2345), .A(n1922), 
        .ZN(n651) );
  AOI22_X2 U1293 ( .A1(n438), .A2(n459), .B1(n439), .B2(n460), .ZN(n1922) );
  OAI221_X2 U1294 ( .B1(n425), .B2(n1855), .C1(n426), .C2(n1850), .A(n1911), 
        .ZN(n1916) );
  OAI221_X2 U1295 ( .B1(n1983), .B2(n2347), .C1(n1991), .C2(n2345), .A(n1923), 
        .ZN(n649) );
  AOI22_X2 U1296 ( .A1(n438), .A2(n463), .B1(n439), .B2(n464), .ZN(n1923) );
  OAI221_X2 U1297 ( .B1(n1989), .B2(n2347), .C1(n1990), .C2(n2344), .A(n1924), 
        .ZN(n1833) );
  AOI22_X2 U1298 ( .A1(n438), .A2(n450), .B1(n439), .B2(n476), .ZN(n1924) );
  OAI221_X2 U1299 ( .B1(n1925), .B2(n719), .C1(n1990), .C2(n634), .A(n1926), 
        .ZN(n1001) );
  AOI22_X2 U1300 ( .A1(sdata[9]), .A2(n2431), .B1(i_dividend[9]), .B2(n2427), 
        .ZN(n1926) );
  OAI22_X2 U1302 ( .A1(n423), .A2(n1869), .B1(n424), .B2(n405), .ZN(n1929) );
  OAI221_X2 U1303 ( .B1(n2005), .B2(n2347), .C1(n2006), .C2(n2344), .A(n1930), 
        .ZN(n661) );
  AOI22_X2 U1304 ( .A1(n438), .A2(n447), .B1(n439), .B2(n452), .ZN(n1930) );
  OAI221_X2 U1305 ( .B1(n2003), .B2(n2347), .C1(n2008), .C2(n2344), .A(n1931), 
        .ZN(n660) );
  AOI22_X2 U1306 ( .A1(n438), .A2(n474), .B1(n439), .B2(n475), .ZN(n1931) );
  OAI22_X2 U1307 ( .A1(n422), .A2(n1907), .B1(n686), .B2(n1908), .ZN(n1928) );
  OAI221_X2 U1309 ( .B1(n1995), .B2(n2347), .C1(n1996), .C2(n2344), .A(n1932), 
        .ZN(n659) );
  AOI22_X2 U1310 ( .A1(n438), .A2(n458), .B1(n439), .B2(n459), .ZN(n1932) );
  OAI221_X2 U1311 ( .B1(n420), .B2(n1855), .C1(n421), .C2(n1850), .A(n1911), 
        .ZN(n1927) );
  OAI221_X2 U1312 ( .B1(n1991), .B2(n2347), .C1(n1992), .C2(n2344), .A(n1933), 
        .ZN(n658) );
  AOI22_X2 U1313 ( .A1(n438), .A2(n462), .B1(n439), .B2(n463), .ZN(n1933) );
  OAI221_X2 U1314 ( .B1(n1990), .B2(n2347), .C1(n1981), .C2(n2344), .A(n1934), 
        .ZN(n1847) );
  AOI22_X2 U1315 ( .A1(n438), .A2(n453), .B1(n439), .B2(n450), .ZN(n1934) );
  OAI221_X2 U1316 ( .B1(n1935), .B2(n719), .C1(n1981), .C2(n2337), .A(n1936), 
        .ZN(n1000) );
  AOI22_X2 U1317 ( .A1(sdata[10]), .A2(n2431), .B1(i_dividend[10]), .B2(n2427), 
        .ZN(n1936) );
  NAND4_X2 U1320 ( .A1(state[1]), .A2(n1651), .A3(n105), .A4(n238), .ZN(n916)
         );
  NAND2_X2 U1323 ( .A1(n106), .A2(n968), .ZN(n719) );
  NAND4_X2 U1325 ( .A1(state[3]), .A2(n1590), .A3(n240), .A4(n2335), .ZN(n963)
         );
  OAI22_X2 U1328 ( .A1(n418), .A2(n1869), .B1(n419), .B2(n405), .ZN(n1939) );
  OAI221_X2 U1330 ( .B1(n2006), .B2(n2347), .C1(n2002), .C2(n2344), .A(n1940), 
        .ZN(n674) );
  AOI22_X2 U1331 ( .A1(n438), .A2(n451), .B1(n439), .B2(n447), .ZN(n1940) );
  NAND2_X2 U1332 ( .A1(n1839), .A2(n404), .ZN(n1869) );
  OAI221_X2 U1334 ( .B1(n2008), .B2(n2347), .C1(n1982), .C2(n2344), .A(n1941), 
        .ZN(n673) );
  AOI22_X2 U1335 ( .A1(n438), .A2(n465), .B1(n439), .B2(n474), .ZN(n1941) );
  OAI22_X2 U1336 ( .A1(n417), .A2(n1907), .B1(n443), .B2(n1908), .ZN(n1938) );
  OR2_X2 U1337 ( .A1(n1836), .A2(n1853), .ZN(n1908) );
  OAI22_X2 U1339 ( .A1(n2000), .A2(n2346), .B1(n870), .B2(n2016), .ZN(n670) );
  NAND2_X2 U1340 ( .A1(n412), .A2(n402), .ZN(n1907) );
  OAI221_X2 U1341 ( .B1(n1996), .B2(n2346), .C1(n1997), .C2(n2344), .A(n1942), 
        .ZN(n671) );
  AOI22_X2 U1342 ( .A1(n438), .A2(n457), .B1(n439), .B2(n458), .ZN(n1942) );
  OAI221_X2 U1343 ( .B1(n415), .B2(n1855), .C1(n416), .C2(n1850), .A(n1911), 
        .ZN(n1937) );
  NAND2_X2 U1345 ( .A1(n401), .A2(n455), .ZN(n1856) );
  NAND2_X2 U1347 ( .A1(n944), .A2(n406), .ZN(n1853) );
  NAND2_X2 U1348 ( .A1(n404), .A2(n1838), .ZN(n1850) );
  OAI221_X2 U1350 ( .B1(n1992), .B2(n2347), .C1(n1993), .C2(n2344), .A(n1943), 
        .ZN(n669) );
  AOI22_X2 U1351 ( .A1(n438), .A2(n461), .B1(n439), .B2(n462), .ZN(n1943) );
  NAND2_X2 U1352 ( .A1(n404), .A2(n412), .ZN(n1855) );
  NAND2_X2 U1354 ( .A1(n945), .A2(n944), .ZN(n718) );
  OAI221_X2 U1355 ( .B1(n1981), .B2(n2346), .C1(n2004), .C2(n2344), .A(n1944), 
        .ZN(n1861) );
  AOI22_X2 U1356 ( .A1(n438), .A2(n449), .B1(n439), .B2(n453), .ZN(n1944) );
  NAND2_X2 U1357 ( .A1(n949), .A2(n441), .ZN(n1843) );
  NAND2_X2 U1358 ( .A1(n445), .A2(n441), .ZN(n1844) );
  INV_X4 U1362 ( .A(n721), .ZN(n4) );
  INV_X4 U1365 ( .A(n1814), .ZN(n7) );
  INV_X4 U1366 ( .A(n1801), .ZN(n8) );
  INV_X4 U1367 ( .A(n1786), .ZN(n9) );
  INV_X4 U1368 ( .A(n1771), .ZN(n10) );
  INV_X4 U1369 ( .A(n1761), .ZN(n11) );
  INV_X4 U1370 ( .A(n1751), .ZN(n12) );
  INV_X4 U1371 ( .A(n1741), .ZN(n13) );
  INV_X4 U1372 ( .A(n1731), .ZN(n14) );
  INV_X4 U1373 ( .A(n1721), .ZN(n15) );
  INV_X4 U1374 ( .A(n1711), .ZN(n16) );
  INV_X4 U1375 ( .A(n1701), .ZN(n17) );
  INV_X4 U1376 ( .A(n1691), .ZN(n18) );
  INV_X4 U1377 ( .A(n1686), .ZN(n19) );
  INV_X4 U1378 ( .A(n1674), .ZN(n20) );
  INV_X4 U1380 ( .A(n762), .ZN(n22) );
  INV_X4 U1381 ( .A(n892), .ZN(n23) );
  INV_X4 U1382 ( .A(n885), .ZN(n24) );
  INV_X4 U1383 ( .A(n878), .ZN(n25) );
  INV_X4 U1384 ( .A(n871), .ZN(n26) );
  INV_X4 U1385 ( .A(n863), .ZN(n27) );
  INV_X4 U1386 ( .A(n837), .ZN(n28) );
  INV_X4 U1387 ( .A(n830), .ZN(n29) );
  INV_X4 U1388 ( .A(n823), .ZN(n30) );
  INV_X4 U1389 ( .A(n816), .ZN(n31) );
  INV_X4 U1390 ( .A(n809), .ZN(n32) );
  INV_X4 U1391 ( .A(n802), .ZN(n33) );
  INV_X4 U1392 ( .A(n795), .ZN(n34) );
  INV_X4 U1393 ( .A(n783), .ZN(n35) );
  INV_X4 U1394 ( .A(n777), .ZN(n36) );
  INV_X4 U1395 ( .A(n899), .ZN(n37) );
  INV_X4 U1399 ( .A(n612), .ZN(n41) );
  INV_X4 U1401 ( .A(n1591), .ZN(n43) );
  INV_X4 U1402 ( .A(n1118), .ZN(n44) );
  INV_X4 U1403 ( .A(n749), .ZN(n45) );
  INV_X4 U1404 ( .A(n747), .ZN(n46) );
  INV_X4 U1405 ( .A(n744), .ZN(n47) );
  INV_X4 U1406 ( .A(n741), .ZN(n48) );
  INV_X4 U1407 ( .A(n738), .ZN(n49) );
  INV_X4 U1408 ( .A(n735), .ZN(n50) );
  INV_X4 U1409 ( .A(n625), .ZN(n51) );
  INV_X4 U1410 ( .A(n623), .ZN(n52) );
  INV_X4 U1411 ( .A(n621), .ZN(n53) );
  INV_X4 U1412 ( .A(n619), .ZN(n54) );
  INV_X4 U1413 ( .A(n617), .ZN(n55) );
  INV_X4 U1414 ( .A(n614), .ZN(n56) );
  INV_X4 U1418 ( .A(n711), .ZN(n60) );
  INV_X4 U1419 ( .A(n678), .ZN(n61) );
  INV_X4 U1421 ( .A(n639), .ZN(n63) );
  INV_X4 U1422 ( .A(n914), .ZN(n64) );
  INV_X4 U1426 ( .A(n610), .ZN(n68) );
  INV_X4 U1427 ( .A(n968), .ZN(n69) );
  INV_X4 U1428 ( .A(n1636), .ZN(n70) );
  INV_X4 U1429 ( .A(n1635), .ZN(n71) );
  INV_X4 U1430 ( .A(n1634), .ZN(n72) );
  INV_X4 U1431 ( .A(n1633), .ZN(n73) );
  INV_X4 U1432 ( .A(n1632), .ZN(n74) );
  INV_X4 U1433 ( .A(n1631), .ZN(n75) );
  INV_X4 U1434 ( .A(n1630), .ZN(n76) );
  INV_X4 U1435 ( .A(n1629), .ZN(n77) );
  INV_X4 U1436 ( .A(n1628), .ZN(n78) );
  INV_X4 U1437 ( .A(n1627), .ZN(n79) );
  INV_X4 U1438 ( .A(n1626), .ZN(n80) );
  INV_X4 U1439 ( .A(n1625), .ZN(n81) );
  INV_X4 U1440 ( .A(n1624), .ZN(n82) );
  INV_X4 U1441 ( .A(n1623), .ZN(n83) );
  INV_X4 U1442 ( .A(n1622), .ZN(n84) );
  INV_X4 U1443 ( .A(n1621), .ZN(n85) );
  INV_X4 U1444 ( .A(n1620), .ZN(n86) );
  INV_X4 U1445 ( .A(n1619), .ZN(n87) );
  INV_X4 U1446 ( .A(n1618), .ZN(n88) );
  INV_X4 U1447 ( .A(n1617), .ZN(n89) );
  INV_X4 U1448 ( .A(n1616), .ZN(n90) );
  INV_X4 U1449 ( .A(n1615), .ZN(n91) );
  INV_X4 U1450 ( .A(n1614), .ZN(n92) );
  INV_X4 U1451 ( .A(n1613), .ZN(n93) );
  INV_X4 U1452 ( .A(n1612), .ZN(n94) );
  INV_X4 U1453 ( .A(n1611), .ZN(n95) );
  INV_X4 U1454 ( .A(n1610), .ZN(n96) );
  INV_X4 U1455 ( .A(n1609), .ZN(n97) );
  INV_X4 U1456 ( .A(n1608), .ZN(n98) );
  INV_X4 U1457 ( .A(n1607), .ZN(n99) );
  INV_X4 U1458 ( .A(n1605), .ZN(n100) );
  INV_X4 U1459 ( .A(n754), .ZN(n101) );
  INV_X4 U1461 ( .A(n913), .ZN(n103) );
  INV_X4 U1462 ( .A(n611), .ZN(n104) );
  INV_X4 U1464 ( .A(n963), .ZN(n106) );
  INV_X4 U1465 ( .A(n964), .ZN(n107) );
  INV_X4 U1478 ( .A(n1650), .ZN(n120) );
  INV_X4 U1528 ( .A(n627), .ZN(o_ready) );
  INV_X4 U1575 ( .A(n1675), .ZN(n217) );
  INV_X4 U1594 ( .A(n593), .ZN(n236) );
  INV_X4 U1600 ( .A(n932), .ZN(n242) );
  INV_X4 U1601 ( .A(n931), .ZN(n243) );
  INV_X4 U1602 ( .A(n920), .ZN(n244) );
  INV_X4 U1603 ( .A(n919), .ZN(n245) );
  INV_X4 U1604 ( .A(n925), .ZN(n246) );
  INV_X4 U1605 ( .A(n924), .ZN(n247) );
  INV_X4 U1606 ( .A(n1445), .ZN(n248) );
  INV_X4 U1607 ( .A(n928), .ZN(n249) );
  INV_X4 U1608 ( .A(n1478), .ZN(n250) );
  INV_X4 U1609 ( .A(n912), .ZN(n251) );
  INV_X4 U1610 ( .A(n907), .ZN(n252) );
  INV_X4 U1611 ( .A(n906), .ZN(n253) );
  INV_X4 U1612 ( .A(n923), .ZN(n254) );
  INV_X4 U1613 ( .A(n909), .ZN(n255) );
  INV_X4 U1614 ( .A(n930), .ZN(n256) );
  INV_X4 U1615 ( .A(n929), .ZN(n257) );
  INV_X4 U1616 ( .A(n908), .ZN(n258) );
  INV_X4 U1617 ( .A(n918), .ZN(n259) );
  INV_X4 U1618 ( .A(n911), .ZN(n260) );
  INV_X4 U1619 ( .A(n910), .ZN(n261) );
  INV_X4 U1620 ( .A(n1466), .ZN(n262) );
  INV_X4 U1621 ( .A(n927), .ZN(n263) );
  INV_X4 U1622 ( .A(n926), .ZN(n264) );
  INV_X4 U1623 ( .A(n922), .ZN(n265) );
  INV_X4 U1624 ( .A(n921), .ZN(n266) );
  INV_X4 U1625 ( .A(n769), .ZN(n267) );
  INV_X4 U1626 ( .A(n905), .ZN(n268) );
  INV_X4 U1627 ( .A(n904), .ZN(n269) );
  INV_X4 U1628 ( .A(n917), .ZN(n270) );
  INV_X4 U1629 ( .A(n1310), .ZN(n271) );
  INV_X4 U1630 ( .A(n1503), .ZN(n272) );
  INV_X4 U1631 ( .A(n1504), .ZN(n273) );
  INV_X4 U1633 ( .A(n903), .ZN(n275) );
  INV_X4 U1634 ( .A(n902), .ZN(n276) );
  INV_X4 U1635 ( .A(n1599), .ZN(n277) );
  INV_X4 U1636 ( .A(n1299), .ZN(n278) );
  INV_X4 U1638 ( .A(n1123), .ZN(n280) );
  INV_X4 U1640 ( .A(n1501), .ZN(n282) );
  INV_X4 U1641 ( .A(n900), .ZN(n283) );
  INV_X4 U1643 ( .A(n729), .ZN(n285) );
  INV_X4 U1644 ( .A(n728), .ZN(n286) );
  INV_X4 U1645 ( .A(n1339), .ZN(n287) );
  INV_X4 U1646 ( .A(n727), .ZN(n288) );
  INV_X4 U1647 ( .A(n726), .ZN(n289) );
  INV_X4 U1648 ( .A(n725), .ZN(n290) );
  INV_X4 U1649 ( .A(n724), .ZN(n291) );
  INV_X4 U1650 ( .A(n723), .ZN(n292) );
  INV_X4 U1651 ( .A(n1341), .ZN(n293) );
  INV_X4 U1652 ( .A(n1324), .ZN(n294) );
  INV_X4 U1653 ( .A(n1359), .ZN(n295) );
  INV_X4 U1654 ( .A(n1334), .ZN(n296) );
  INV_X4 U1655 ( .A(n1307), .ZN(n297) );
  INV_X4 U1657 ( .A(n737), .ZN(n299) );
  INV_X4 U1658 ( .A(n1394), .ZN(n300) );
  INV_X4 U1659 ( .A(n734), .ZN(n301) );
  INV_X4 U1660 ( .A(n733), .ZN(n302) );
  INV_X4 U1661 ( .A(n1371), .ZN(n303) );
  INV_X4 U1662 ( .A(n732), .ZN(n304) );
  INV_X4 U1663 ( .A(n731), .ZN(n305) );
  INV_X4 U1664 ( .A(n1363), .ZN(n306) );
  INV_X4 U1665 ( .A(n730), .ZN(n307) );
  INV_X4 U1666 ( .A(n1427), .ZN(n308) );
  INV_X4 U1667 ( .A(n1357), .ZN(n309) );
  INV_X4 U1668 ( .A(n1413), .ZN(n310) );
  INV_X4 U1669 ( .A(n1377), .ZN(n311) );
  INV_X4 U1670 ( .A(n1351), .ZN(n312) );
  INV_X4 U1671 ( .A(n1407), .ZN(n313) );
  INV_X4 U1672 ( .A(n740), .ZN(n314) );
  INV_X4 U1673 ( .A(n1415), .ZN(n315) );
  INV_X4 U1674 ( .A(n1434), .ZN(n316) );
  INV_X4 U1675 ( .A(n743), .ZN(n317) );
  INV_X4 U1676 ( .A(n1436), .ZN(n318) );
  INV_X4 U1677 ( .A(n1454), .ZN(n319) );
  INV_X4 U1678 ( .A(n1429), .ZN(n320) );
  INV_X4 U1679 ( .A(n1447), .ZN(n321) );
  INV_X4 U1681 ( .A(n746), .ZN(n323) );
  INV_X4 U1682 ( .A(n1456), .ZN(n324) );
  INV_X4 U1683 ( .A(n1483), .ZN(n325) );
  INV_X4 U1684 ( .A(n1449), .ZN(n326) );
  INV_X4 U1685 ( .A(n1474), .ZN(n327) );
  INV_X4 U1686 ( .A(n1482), .ZN(n328) );
  INV_X4 U1687 ( .A(n1510), .ZN(n329) );
  INV_X4 U1688 ( .A(n751), .ZN(n330) );
  INV_X4 U1689 ( .A(n1517), .ZN(n331) );
  INV_X4 U1690 ( .A(n1507), .ZN(n332) );
  INV_X4 U1691 ( .A(n1485), .ZN(n333) );
  INV_X4 U1692 ( .A(n1476), .ZN(n334) );
  INV_X4 U1698 ( .A(n1346), .ZN(n340) );
  INV_X4 U1699 ( .A(n1396), .ZN(n341) );
  INV_X4 U1701 ( .A(n1331), .ZN(n343) );
  INV_X4 U1702 ( .A(n1365), .ZN(n344) );
  INV_X4 U1704 ( .A(n753), .ZN(n346) );
  INV_X4 U1705 ( .A(n752), .ZN(n347) );
  INV_X4 U1706 ( .A(n1580), .ZN(n348) );
  INV_X4 U1707 ( .A(n1555), .ZN(n349) );
  INV_X4 U1708 ( .A(n1516), .ZN(n350) );
  INV_X4 U1709 ( .A(n1588), .ZN(n351) );
  INV_X4 U1711 ( .A(n1509), .ZN(n353) );
  INV_X4 U1712 ( .A(n1512), .ZN(n354) );
  INV_X4 U1713 ( .A(n1389), .ZN(n355) );
  INV_X4 U1714 ( .A(n1332), .ZN(n356) );
  INV_X4 U1715 ( .A(n1379), .ZN(n357) );
  INV_X4 U1716 ( .A(n1373), .ZN(n358) );
  INV_X4 U1722 ( .A(n1552), .ZN(n364) );
  INV_X4 U1724 ( .A(n1120), .ZN(n366) );
  INV_X4 U1725 ( .A(n1117), .ZN(n367) );
  INV_X4 U1726 ( .A(n1586), .ZN(n368) );
  INV_X4 U1727 ( .A(n1576), .ZN(n369) );
  INV_X4 U1729 ( .A(n1581), .ZN(n371) );
  INV_X4 U1758 ( .A(n1856), .ZN(n400) );
  INV_X4 U1760 ( .A(n1853), .ZN(n402) );
  INV_X4 U1761 ( .A(n1869), .ZN(n403) );
  INV_X4 U1762 ( .A(n718), .ZN(n404) );
  INV_X4 U1763 ( .A(n1872), .ZN(n405) );
  INV_X4 U1765 ( .A(n702), .ZN(n407) );
  INV_X4 U1766 ( .A(n700), .ZN(n408) );
  INV_X4 U1767 ( .A(n698), .ZN(n409) );
  INV_X4 U1768 ( .A(n1878), .ZN(n410) );
  INV_X4 U1769 ( .A(n682), .ZN(n411) );
  INV_X4 U1770 ( .A(n672), .ZN(n412) );
  INV_X4 U1771 ( .A(n667), .ZN(n413) );
  INV_X4 U1773 ( .A(n1861), .ZN(n415) );
  INV_X4 U1774 ( .A(n669), .ZN(n416) );
  INV_X4 U1775 ( .A(n671), .ZN(n417) );
  INV_X4 U1776 ( .A(n673), .ZN(n418) );
  INV_X4 U1777 ( .A(n674), .ZN(n419) );
  INV_X4 U1778 ( .A(n1847), .ZN(n420) );
  INV_X4 U1779 ( .A(n658), .ZN(n421) );
  INV_X4 U1780 ( .A(n659), .ZN(n422) );
  INV_X4 U1781 ( .A(n660), .ZN(n423) );
  INV_X4 U1782 ( .A(n661), .ZN(n424) );
  INV_X4 U1783 ( .A(n1833), .ZN(n425) );
  INV_X4 U1784 ( .A(n649), .ZN(n426) );
  INV_X4 U1785 ( .A(n651), .ZN(n427) );
  INV_X4 U1786 ( .A(n650), .ZN(n428) );
  INV_X4 U1787 ( .A(n652), .ZN(n429) );
  INV_X4 U1788 ( .A(n653), .ZN(n430) );
  INV_X4 U1789 ( .A(n1873), .ZN(n431) );
  INV_X4 U1790 ( .A(n636), .ZN(n432) );
  INV_X4 U1791 ( .A(n640), .ZN(n433) );
  INV_X4 U1792 ( .A(n638), .ZN(n434) );
  INV_X4 U1793 ( .A(n642), .ZN(n435) );
  INV_X4 U1794 ( .A(n644), .ZN(n436) );
  INV_X4 U1795 ( .A(n1834), .ZN(n437) );
  INV_X4 U1798 ( .A(n686), .ZN(n440) );
  INV_X4 U1801 ( .A(n670), .ZN(n443) );
  INV_X4 U1839 ( .A(n1506), .ZN(n481) );
  INV_X4 U1840 ( .A(n1350), .ZN(n482) );
  INV_X4 U1843 ( .A(n1538), .ZN(n485) );
  INV_X4 U1848 ( .A(n1355), .ZN(n490) );
  INV_X4 U1852 ( .A(n1541), .ZN(n494) );
  INV_X4 U1853 ( .A(n1564), .ZN(n495) );
  INV_X4 U1854 ( .A(n1535), .ZN(n496) );
  INV_X4 U1856 ( .A(n1369), .ZN(n498) );
  INV_X4 U1859 ( .A(n1461), .ZN(n501) );
  INV_X4 U1861 ( .A(n954), .ZN(n503) );
  INV_X4 U1862 ( .A(n1532), .ZN(n504) );
  INV_X4 U1864 ( .A(n1530), .ZN(n506) );
  INV_X4 U1865 ( .A(n1401), .ZN(n507) );
  INV_X4 U1866 ( .A(n1444), .ZN(n508) );
  INV_X4 U1867 ( .A(n1393), .ZN(n509) );
  INV_X4 U1870 ( .A(n1529), .ZN(n512) );
  INV_X4 U1873 ( .A(n1495), .ZN(n515) );
  INV_X4 U1874 ( .A(n1527), .ZN(n516) );
  INV_X4 U1878 ( .A(n1544), .ZN(n520) );
  INV_X4 U1879 ( .A(n956), .ZN(n521) );
  INV_X4 U1881 ( .A(n1542), .ZN(n523) );
  INV_X4 U1885 ( .A(n952), .ZN(n527) );
  INV_X4 U1886 ( .A(n960), .ZN(n528) );
  INV_X4 U1888 ( .A(n953), .ZN(n530) );
  INV_X4 U1897 ( .A(i_dividend[31]), .ZN(n539) );
  INV_X4 U1898 ( .A(i_dividend[30]), .ZN(n540) );
  INV_X4 U1899 ( .A(i_dividend[29]), .ZN(n541) );
  INV_X4 U1900 ( .A(i_dividend[28]), .ZN(n542) );
  INV_X4 U1901 ( .A(i_dividend[27]), .ZN(n543) );
  INV_X4 U1902 ( .A(i_dividend[22]), .ZN(n544) );
  INV_X4 U1903 ( .A(i_dividend[21]), .ZN(n545) );
  INV_X4 U1904 ( .A(i_dividend[20]), .ZN(n546) );
  INV_X4 U1905 ( .A(i_dividend[18]), .ZN(n547) );
  INV_X4 U1906 ( .A(i_dividend[16]), .ZN(n548) );
  INV_X4 U1907 ( .A(i_divisor[31]), .ZN(n549) );
  INV_X4 U1908 ( .A(i_divisor[30]), .ZN(n550) );
  INV_X4 U1909 ( .A(i_divisor[29]), .ZN(n551) );
  INV_X4 U1910 ( .A(i_divisor[28]), .ZN(n552) );
  INV_X4 U1911 ( .A(i_divisor[27]), .ZN(n553) );
  INV_X4 U1912 ( .A(i_divisor[26]), .ZN(n554) );
  INV_X4 U1913 ( .A(i_divisor[25]), .ZN(n555) );
  INV_X4 U1914 ( .A(i_divisor[24]), .ZN(n556) );
  INV_X4 U1915 ( .A(i_divisor[23]), .ZN(n557) );
  INV_X4 U1916 ( .A(i_divisor[22]), .ZN(n558) );
  INV_X4 U1917 ( .A(i_divisor[21]), .ZN(n559) );
  INV_X4 U1918 ( .A(i_divisor[20]), .ZN(n560) );
  INV_X4 U1919 ( .A(i_divisor[19]), .ZN(n561) );
  INV_X4 U1920 ( .A(i_divisor[18]), .ZN(n562) );
  INV_X4 U1921 ( .A(i_divisor[17]), .ZN(n563) );
  INV_X4 U1922 ( .A(i_divisor[16]), .ZN(n564) );
  INV_X4 U1923 ( .A(i_divisor[15]), .ZN(n565) );
  INV_X4 U1924 ( .A(i_divisor[14]), .ZN(n566) );
  INV_X4 U1925 ( .A(i_divisor[13]), .ZN(n567) );
  INV_X4 U1926 ( .A(i_divisor[12]), .ZN(n568) );
  INV_X4 U1927 ( .A(i_divisor[11]), .ZN(n569) );
  INV_X4 U1928 ( .A(i_divisor[10]), .ZN(n570) );
  INV_X4 U1929 ( .A(i_divisor[9]), .ZN(n571) );
  INV_X4 U1930 ( .A(i_divisor[8]), .ZN(n572) );
  INV_X4 U1931 ( .A(i_divisor[7]), .ZN(n573) );
  INV_X4 U1932 ( .A(i_divisor[6]), .ZN(n574) );
  INV_X4 U1933 ( .A(i_divisor[5]), .ZN(n575) );
  INV_X4 U1934 ( .A(i_divisor[4]), .ZN(n576) );
  INV_X4 U1935 ( .A(i_divisor[3]), .ZN(n577) );
  INV_X4 U1936 ( .A(i_divisor[2]), .ZN(n578) );
  INV_X4 U1937 ( .A(i_divisor[1]), .ZN(n579) );
  INV_X4 U1938 ( .A(i_divisor[0]), .ZN(n580) );
  OAI33_X1 U1939 ( .A1(n1558), .A2(n1362), .A3(n1441), .B1(n528), .B2(n515), 
        .B3(n523), .ZN(n1560) );
  SDFFR_X2 o_remainder_reg_1_ ( .D(n1261), .SI(o_remainder[0]), .SE(test_se), 
        .CK(i_clk), .RN(n2451), .Q(o_remainder[1]), .QN(n2638) );
  SDFFR_X2 o_remainder_reg_0_ ( .D(n1262), .SI(o_quotient[31]), .SE(test_se), 
        .CK(i_clk), .RN(n2445), .Q(o_remainder[0]), .QN(n2637) );
  SDFFR_X2 o_remainder_reg_2_ ( .D(n1260), .SI(o_remainder[1]), .SE(test_se), 
        .CK(i_clk), .RN(n2445), .Q(o_remainder[2]), .QN(n2639) );
  SDFFR_X2 o_quotient_reg_2_ ( .D(n1222), .SI(o_quotient[1]), .SE(test_se), 
        .CK(i_clk), .RN(n2445), .Q(o_quotient[2]), .QN(n2671) );
  SDFFR_X2 o_quotient_reg_1_ ( .D(n1223), .SI(o_quotient[0]), .SE(test_se), 
        .CK(i_clk), .RN(n2445), .Q(o_quotient[1]), .QN(n2670) );
  SDFFR_X2 o_quotient_reg_0_ ( .D(n1224), .SI(nq[30]), .SE(test_se), .CK(i_clk), .RN(n2445), .Q(o_quotient[0]), .QN(n2669) );
  SDFFR_X2 o_quotient_reg_3_ ( .D(n1221), .SI(o_quotient[2]), .SE(test_se), 
        .CK(i_clk), .RN(n2445), .Q(o_quotient[3]), .QN(n2672) );
  SDFFR_X2 o_remainder_reg_3_ ( .D(n1259), .SI(o_remainder[2]), .SE(test_se), 
        .CK(i_clk), .RN(n2445), .Q(o_remainder[3]), .QN(n2640) );
  SDFFR_X2 o_quotient_reg_5_ ( .D(n1219), .SI(o_quotient[4]), .SE(test_se), 
        .CK(i_clk), .RN(n2445), .Q(o_quotient[5]), .QN(n2674) );
  SDFFR_X2 o_remainder_reg_5_ ( .D(n1257), .SI(o_remainder[4]), .SE(test_se), 
        .CK(i_clk), .RN(n2446), .Q(o_remainder[5]), .QN(n2642) );
  SDFFR_X2 o_quotient_reg_4_ ( .D(n1220), .SI(o_quotient[3]), .SE(test_se), 
        .CK(i_clk), .RN(n2446), .Q(o_quotient[4]), .QN(n2673) );
  SDFFR_X2 o_remainder_reg_4_ ( .D(n1258), .SI(o_remainder[3]), .SE(test_se), 
        .CK(i_clk), .RN(n2446), .Q(o_remainder[4]), .QN(n2641) );
  SDFFR_X2 o_quotient_reg_7_ ( .D(n1217), .SI(o_quotient[6]), .SE(test_se), 
        .CK(i_clk), .RN(n2446), .Q(o_quotient[7]), .QN(n2676) );
  SDFFR_X2 o_remainder_reg_7_ ( .D(n1255), .SI(o_remainder[6]), .SE(test_se), 
        .CK(i_clk), .RN(n2446), .Q(o_remainder[7]), .QN(n2644) );
  SDFFR_X2 o_quotient_reg_6_ ( .D(n1218), .SI(o_quotient[5]), .SE(test_se), 
        .CK(i_clk), .RN(n2447), .Q(o_quotient[6]), .QN(n2675) );
  SDFFR_X2 o_remainder_reg_6_ ( .D(n1256), .SI(o_remainder[5]), .SE(test_se), 
        .CK(i_clk), .RN(n2447), .Q(o_remainder[6]), .QN(n2643) );
  SDFFR_X2 o_quotient_reg_13_ ( .D(n1211), .SI(o_quotient[12]), .SE(test_se), 
        .CK(i_clk), .RN(n2447), .Q(o_quotient[13]), .QN(n2682) );
  SDFFR_X2 o_quotient_reg_11_ ( .D(n1213), .SI(o_quotient[10]), .SE(test_se), 
        .CK(i_clk), .RN(n2447), .Q(o_quotient[11]), .QN(n2680) );
  SDFFR_X2 o_quotient_reg_9_ ( .D(n1215), .SI(o_quotient[8]), .SE(test_se), 
        .CK(i_clk), .RN(n2447), .Q(o_quotient[9]), .QN(n2678) );
  SDFFR_X2 o_remainder_reg_13_ ( .D(n1249), .SI(o_remainder[12]), .SE(test_se), 
        .CK(i_clk), .RN(n2447), .Q(o_remainder[13]), .QN(n2650) );
  SDFFR_X2 o_remainder_reg_11_ ( .D(n1251), .SI(o_remainder[10]), .SE(test_se), 
        .CK(i_clk), .RN(n2447), .Q(o_remainder[11]), .QN(n2648) );
  SDFFR_X2 o_remainder_reg_9_ ( .D(n1253), .SI(o_remainder[8]), .SE(test_se), 
        .CK(i_clk), .RN(n2447), .Q(o_remainder[9]), .QN(n2646) );
  SDFFR_X2 o_quotient_reg_8_ ( .D(n1216), .SI(o_quotient[7]), .SE(test_se), 
        .CK(i_clk), .RN(n2448), .Q(o_quotient[8]), .QN(n2677) );
  SDFFR_X2 o_remainder_reg_8_ ( .D(n1254), .SI(o_remainder[7]), .SE(test_se), 
        .CK(i_clk), .RN(n2448), .Q(o_remainder[8]), .QN(n2645) );
  SDFFR_X2 o_quotient_reg_15_ ( .D(n1209), .SI(o_quotient[14]), .SE(test_se), 
        .CK(i_clk), .RN(n2450), .Q(o_quotient[15]), .QN(n2684) );
  SDFFR_X2 o_remainder_reg_15_ ( .D(n1247), .SI(o_remainder[14]), .SE(test_se), 
        .CK(i_clk), .RN(n2450), .Q(o_remainder[15]), .QN(n2652) );
  SDFFR_X2 o_quotient_reg_14_ ( .D(n1210), .SI(o_quotient[13]), .SE(test_se), 
        .CK(i_clk), .RN(n2450), .Q(o_quotient[14]), .QN(n2683) );
  SDFFR_X2 o_quotient_reg_12_ ( .D(n1212), .SI(o_quotient[11]), .SE(test_se), 
        .CK(i_clk), .RN(n2450), .Q(o_quotient[12]), .QN(n2681) );
  SDFFR_X2 o_quotient_reg_10_ ( .D(n1214), .SI(o_quotient[9]), .SE(test_se), 
        .CK(i_clk), .RN(n2450), .Q(o_quotient[10]), .QN(n2679) );
  SDFFR_X2 o_remainder_reg_14_ ( .D(n1248), .SI(o_remainder[13]), .SE(test_se), 
        .CK(i_clk), .RN(n2450), .Q(o_remainder[14]), .QN(n2651) );
  SDFFR_X2 o_remainder_reg_12_ ( .D(n1250), .SI(o_remainder[11]), .SE(test_se), 
        .CK(i_clk), .RN(n2450), .Q(o_remainder[12]), .QN(n2649) );
  SDFFR_X2 o_remainder_reg_10_ ( .D(n1252), .SI(o_remainder[9]), .SE(test_se), 
        .CK(i_clk), .RN(n2450), .Q(o_remainder[10]), .QN(n2647) );
  SDFFR_X2 o_quotient_reg_16_ ( .D(n1208), .SI(o_quotient[15]), .SE(test_se), 
        .CK(i_clk), .RN(n2450), .Q(o_quotient[16]), .QN(n2685) );
  SDFFR_X2 o_remainder_reg_16_ ( .D(n1246), .SI(o_remainder[15]), .SE(test_se), 
        .CK(i_clk), .RN(n2451), .Q(o_remainder[16]), .QN(n2653) );
  SDFFR_X2 o_quotient_reg_23_ ( .D(n1201), .SI(o_quotient[22]), .SE(test_se), 
        .CK(i_clk), .RN(n2451), .Q(o_quotient[23]), .QN(n2692) );
  SDFFR_X2 o_quotient_reg_21_ ( .D(n1203), .SI(o_quotient[20]), .SE(test_se), 
        .CK(i_clk), .RN(n2451), .Q(o_quotient[21]), .QN(n2690) );
  SDFFR_X2 o_quotient_reg_19_ ( .D(n1205), .SI(o_quotient[18]), .SE(test_se), 
        .CK(i_clk), .RN(n2451), .Q(o_quotient[19]), .QN(n2688) );
  SDFFR_X2 o_quotient_reg_17_ ( .D(n1207), .SI(o_quotient[16]), .SE(test_se), 
        .CK(i_clk), .RN(n2451), .Q(o_quotient[17]), .QN(n2686) );
  SDFFR_X2 o_remainder_reg_23_ ( .D(n1239), .SI(o_remainder[22]), .SE(test_se), 
        .CK(i_clk), .RN(n2451), .Q(o_remainder[23]), .QN(n2660) );
  SDFFR_X2 o_remainder_reg_21_ ( .D(n1241), .SI(o_remainder[20]), .SE(test_se), 
        .CK(i_clk), .RN(n2451), .Q(o_remainder[21]), .QN(n2658) );
  SDFFR_X2 o_remainder_reg_19_ ( .D(n1243), .SI(o_remainder[18]), .SE(test_se), 
        .CK(i_clk), .RN(n2451), .Q(o_remainder[19]), .QN(n2656) );
  SDFFR_X2 o_remainder_reg_17_ ( .D(n1245), .SI(o_remainder[16]), .SE(test_se), 
        .CK(i_clk), .RN(n2451), .Q(o_remainder[17]), .QN(n2654) );
  SDFFR_X2 o_quotient_reg_27_ ( .D(n1197), .SI(o_quotient[26]), .SE(test_se), 
        .CK(i_clk), .RN(n2452), .Q(o_quotient[27]), .QN(n2696) );
  SDFFR_X2 o_quotient_reg_25_ ( .D(n1199), .SI(o_quotient[24]), .SE(test_se), 
        .CK(i_clk), .RN(n2452), .Q(o_quotient[25]), .QN(n2694) );
  SDFFR_X2 o_remainder_reg_27_ ( .D(n1235), .SI(o_remainder[26]), .SE(test_se), 
        .CK(i_clk), .RN(n2452), .Q(o_remainder[27]), .QN(n2664) );
  SDFFR_X2 o_remainder_reg_25_ ( .D(n1237), .SI(o_remainder[24]), .SE(test_se), 
        .CK(i_clk), .RN(n2452), .Q(o_remainder[25]), .QN(n2662) );
  SDFFR_X2 o_remainder_reg_31_ ( .D(n1231), .SI(q[27]), .SE(test_se), .CK(
        i_clk), .RN(n2452), .Q(o_remainder[31]), .QN(n2668) );
  SDFFR_X2 o_quotient_reg_29_ ( .D(n1195), .SI(o_quotient[28]), .SE(test_se), 
        .CK(i_clk), .RN(n2452), .Q(o_quotient[29]), .QN(n2698) );
  SDFFR_X2 o_remainder_reg_29_ ( .D(n1233), .SI(o_remainder[28]), .SE(test_se), 
        .CK(i_clk), .RN(n2452), .Q(o_remainder[29]), .QN(n2666) );
  SDFFR_X2 o_quotient_reg_31_ ( .D(n1193), .SI(o_quotient[30]), .SE(test_se), 
        .CK(i_clk), .RN(n2452), .Q(o_quotient[31]), .QN(n2700) );
  SDFFR_X2 o_quotient_reg_24_ ( .D(n1200), .SI(o_quotient[23]), .SE(test_se), 
        .CK(i_clk), .RN(n2452), .Q(o_quotient[24]), .QN(n2693) );
  SDFFR_X2 o_quotient_reg_22_ ( .D(n1202), .SI(o_quotient[21]), .SE(test_se), 
        .CK(i_clk), .RN(n2452), .Q(o_quotient[22]), .QN(n2691) );
  SDFFR_X2 o_quotient_reg_20_ ( .D(n1204), .SI(o_quotient[19]), .SE(test_se), 
        .CK(i_clk), .RN(n2452), .Q(o_quotient[20]), .QN(n2689) );
  SDFFR_X2 o_quotient_reg_18_ ( .D(n1206), .SI(o_quotient[17]), .SE(test_se), 
        .CK(i_clk), .RN(n2453), .Q(o_quotient[18]), .QN(n2687) );
  SDFFR_X2 o_remainder_reg_24_ ( .D(n1238), .SI(o_remainder[23]), .SE(test_se), 
        .CK(i_clk), .RN(n2453), .Q(o_remainder[24]), .QN(n2661) );
  SDFFR_X2 o_remainder_reg_22_ ( .D(n1240), .SI(o_remainder[21]), .SE(test_se), 
        .CK(i_clk), .RN(n2453), .Q(o_remainder[22]), .QN(n2659) );
  SDFFR_X2 o_remainder_reg_20_ ( .D(n1242), .SI(o_remainder[19]), .SE(test_se), 
        .CK(i_clk), .RN(n2453), .Q(o_remainder[20]), .QN(n2657) );
  SDFFR_X2 o_remainder_reg_18_ ( .D(n1244), .SI(o_remainder[17]), .SE(test_se), 
        .CK(i_clk), .RN(n2453), .Q(o_remainder[18]), .QN(n2655) );
  SDFFR_X2 o_quotient_reg_28_ ( .D(n1196), .SI(o_quotient[27]), .SE(test_se), 
        .CK(i_clk), .RN(n2453), .Q(o_quotient[28]), .QN(n2697) );
  SDFFR_X2 o_quotient_reg_26_ ( .D(n1198), .SI(o_quotient[25]), .SE(test_se), 
        .CK(i_clk), .RN(n2453), .Q(o_quotient[26]), .QN(n2695) );
  SDFFR_X2 o_remainder_reg_28_ ( .D(n1234), .SI(o_remainder[27]), .SE(test_se), 
        .CK(i_clk), .RN(n2453), .Q(o_remainder[28]), .QN(n2665) );
  SDFFR_X2 o_remainder_reg_26_ ( .D(n1236), .SI(o_remainder[25]), .SE(test_se), 
        .CK(i_clk), .RN(n2453), .Q(o_remainder[26]), .QN(n2663) );
  SDFFR_X2 o_quotient_reg_30_ ( .D(n1194), .SI(o_quotient[29]), .SE(test_se), 
        .CK(i_clk), .RN(n2454), .Q(o_quotient[30]), .QN(n2699) );
  SDFFR_X2 o_remainder_reg_30_ ( .D(n1232), .SI(o_remainder[29]), .SE(test_se), 
        .CK(i_clk), .RN(n2454), .Q(o_remainder[30]), .QN(n2667) );
  SDFFS_X1 state_reg_0_ ( .D(n1191), .SI(n2957), .SE(test_se), .CK(i_clk), 
        .SN(i_rst), .Q(state[0]), .QN(n105) );
  SDFFR_X2 PR_reg_31_ ( .D(n2015), .SI(n154), .SE(test_se), .CK(i_clk), .RN(
        i_rst), .Q(n284), .QN(n3185) );
  SDFFR_X2 ct_reg_2_ ( .D(n2012), .SI(n393), .SE(test_se), .CK(i_clk), .RN(
        n2445), .Q(n396), .QN(n937) );
  SDFFR_X2 ct_reg_1_ ( .D(n2009), .SI(n939), .SE(test_se), .CK(i_clk), .RN(
        n2445), .Q(n393), .QN(n938) );
  SDFFR_X2 ct_reg_0_ ( .D(n2010), .SI(n401), .SE(test_se), .CK(i_clk), .RN(
        n2445), .Q(n394), .QN(n939) );
  SDFFR_X2 ct_reg_3_ ( .D(n2013), .SI(n396), .SE(test_se), .CK(i_clk), .RN(
        n2446), .Q(n397), .QN(n936) );
  SDFFR_X2 ct_reg_5_ ( .D(n2014), .SI(n454), .SE(test_se), .CK(i_clk), .RN(
        n2450), .Q(n479), .QN(n934) );
  SDFFR_X2 ct_reg_4_ ( .D(n2011), .SI(n397), .SE(test_se), .CK(i_clk), .RN(
        n2448), .Q(n454), .QN(n935) );
  SDFFR_X2 ct_1_reg_5_ ( .D(n1106), .SI(n406), .SE(test_se), .CK(i_clk), .RN(
        n2446), .Q(n401), .QN(n944) );
  SDFFR_X2 ct_1_reg_4_ ( .D(n1107), .SI(n3000), .SE(test_se), .CK(i_clk), .RN(
        n2446), .Q(n406), .QN(n945) );
  SDFFR_X2 ct_1_reg_3_ ( .D(n1108), .SI(n414), .SE(test_se), .CK(i_clk), .RN(
        n2446), .Q(n3000), .QN(n946) );
  SDFFR_X2 ct_1_reg_2_ ( .D(n1109), .SI(n948), .SE(test_se), .CK(i_clk), .RN(
        n2446), .Q(n414), .QN(n947) );
  SDFFR_X2 ct_1_reg_1_ ( .D(n1110), .SI(n445), .SE(test_se), .CK(i_clk), .RN(
        n2446), .Q(n441), .QN(n948) );
  SDFFR_X2 ct_1_reg_0_ ( .D(n1111), .SI(n1976), .SE(test_se), .CK(i_clk), .RN(
        n2447), .Q(n445), .QN(n949) );
  SDFFR_X2 nq_reg_1_ ( .D(n1104), .SI(n399), .SE(test_se), .CK(i_clk), .RN(
        n2446), .Q(n2999), .QN(n3284) );
  SDFFR_X2 nq_reg_0_ ( .D(n1105), .SI(n479), .SE(test_se), .CK(i_clk), .RN(
        n2446), .Q(n399), .QN(n3285) );
  SDFFR_X2 PR_1_reg_10_ ( .D(n1000), .SI(n467), .SE(test_se), .CK(i_clk), .RN(
        n2450), .Q(n476), .QN(n1981) );
  SDFFR_X2 PR_1_reg_9_ ( .D(n1001), .SI(n468), .SE(test_se), .CK(i_clk), .RN(
        n2449), .Q(n467), .QN(n1990) );
  SDFFR_X2 PR_1_reg_8_ ( .D(n1002), .SI(n469), .SE(test_se), .CK(i_clk), .RN(
        n2449), .Q(n468), .QN(n1989) );
  SDFFR_X2 PR_1_reg_7_ ( .D(n1003), .SI(n470), .SE(test_se), .CK(i_clk), .RN(
        n2449), .Q(n469), .QN(n1988) );
  SDFFR_X2 shifted_reg_3_ ( .D(n1187), .SI(n2958), .SE(test_se), .CK(i_clk), 
        .RN(n2467), .Q(n2957), .QN(n3119) );
  SDFFR_X2 PR_1_reg_31_ ( .D(n979), .SI(n2000), .SE(test_se), .CK(i_clk), .RN(
        n2448), .Q(n455), .QN(n870) );
  SDFFR_X2 PR_1_reg_14_ ( .D(n996), .SI(n449), .SE(test_se), .CK(i_clk), .RN(
        n2447), .Q(n448), .QN(n2006) );
  SDFFR_X2 PR_1_reg_11_ ( .D(n999), .SI(n476), .SE(test_se), .CK(i_clk), .RN(
        n2448), .Q(n450), .QN(n2004) );
  SDFFR_X2 PR_1_reg_13_ ( .D(n997), .SI(n453), .SE(test_se), .CK(i_clk), .RN(
        n2447), .Q(n449), .QN(n2005) );
  SDFFR_X2 PR_1_reg_12_ ( .D(n998), .SI(n450), .SE(test_se), .CK(i_clk), .RN(
        n2448), .Q(n453), .QN(n2001) );
  SDFFR_X2 PR_1_reg_18_ ( .D(n992), .SI(n451), .SE(test_se), .CK(i_clk), .RN(
        n2447), .Q(n446), .QN(n2008) );
  SDFFR_X2 shifted_reg_2_ ( .D(n1188), .SI(n2959), .SE(test_se), .CK(i_clk), 
        .RN(n2467), .Q(n2958), .QN(n3118) );
  SDFFR_X2 shifted_reg_1_ ( .D(n1189), .SI(n2960), .SE(test_se), .CK(i_clk), 
        .RN(n2467), .Q(n2959), .QN(n3117) );
  SDFFR_X2 PR_1_reg_22_ ( .D(n988), .SI(n465), .SE(test_se), .CK(i_clk), .RN(
        n2449), .Q(n464), .QN(n1992) );
  SDFFR_X2 PR_1_reg_21_ ( .D(n989), .SI(n1983), .SE(test_se), .CK(i_clk), .RN(
        n2449), .Q(n465), .QN(n1991) );
  SDFFR_X2 PR_1_reg_20_ ( .D(n990), .SI(n1982), .SE(test_se), .CK(i_clk), .RN(
        n2449), .Q(n474), .QN(n1983) );
  SDFFR_X2 PR_1_reg_16_ ( .D(n994), .SI(n452), .SE(test_se), .CK(i_clk), .RN(
        n2447), .Q(n447), .QN(n2007) );
  SDFFR_X2 PR_1_reg_19_ ( .D(n991), .SI(n446), .SE(test_se), .CK(i_clk), .RN(
        n2449), .Q(n475), .QN(n1982) );
  SDFFR_X2 PR_1_reg_17_ ( .D(n993), .SI(n447), .SE(test_se), .CK(i_clk), .RN(
        n2448), .Q(n451), .QN(n2003) );
  SDFFR_X2 PR_1_reg_4_ ( .D(n1006), .SI(n477), .SE(test_se), .CK(i_clk), .RN(
        n2449), .Q(n472), .QN(n1985) );
  SDFFR_X2 PR_1_reg_15_ ( .D(n995), .SI(n448), .SE(test_se), .CK(i_clk), .RN(
        n2448), .Q(n452), .QN(n2002) );
  SDFFR_X2 PR_1_reg_0_ ( .D(n1010), .SI(n119), .SE(test_se), .CK(i_clk), .RN(
        n2449), .Q(n466), .QN(n1978) );
  SDFFR_X2 PR_1_reg_6_ ( .D(n1004), .SI(n471), .SE(test_se), .CK(i_clk), .RN(
        n2449), .Q(n470), .QN(n1987) );
  SDFFR_X2 PR_1_reg_5_ ( .D(n1005), .SI(n472), .SE(test_se), .CK(i_clk), .RN(
        n2449), .Q(n471), .QN(n1986) );
  SDFFR_X2 PR_1_reg_29_ ( .D(n981), .SI(n458), .SE(test_se), .CK(i_clk), .RN(
        n2448), .Q(n457), .QN(n1999) );
  SDFFR_X2 PR_1_reg_27_ ( .D(n983), .SI(n460), .SE(test_se), .CK(i_clk), .RN(
        n2448), .Q(n459), .QN(n1997) );
  SDFFR_X2 PR_1_reg_30_ ( .D(n980), .SI(n1999), .SE(test_se), .CK(i_clk), .RN(
        n2448), .Q(n456), .QN(n2000) );
  SDFFR_X2 PR_1_reg_24_ ( .D(n986), .SI(n463), .SE(test_se), .CK(i_clk), .RN(
        n2449), .Q(n462), .QN(n1994) );
  SDFFR_X2 PR_1_reg_26_ ( .D(n984), .SI(n461), .SE(test_se), .CK(i_clk), .RN(
        n2448), .Q(n460), .QN(n1996) );
  SDFFR_X2 PR_1_reg_23_ ( .D(n987), .SI(n464), .SE(test_se), .CK(i_clk), .RN(
        n2449), .Q(n463), .QN(n1993) );
  SDFFR_X2 PR_1_reg_25_ ( .D(n985), .SI(n462), .SE(test_se), .CK(i_clk), .RN(
        n2448), .Q(n461), .QN(n1995) );
  SDFFR_X2 PR_1_reg_28_ ( .D(n982), .SI(n459), .SE(test_se), .CK(i_clk), .RN(
        n2448), .Q(n458), .QN(n1998) );
  SDFFR_X2 PR_1_reg_1_ ( .D(n1009), .SI(n1978), .SE(test_se), .CK(i_clk), .RN(
        n2450), .Q(n478), .QN(n1979) );
  SDFFR_X2 PR_1_reg_2_ ( .D(n1008), .SI(n1979), .SE(test_se), .CK(i_clk), .RN(
        n2449), .Q(n473), .QN(n1984) );
  SDFFR_X2 PR_1_reg_3_ ( .D(n1007), .SI(n473), .SE(test_se), .CK(i_clk), .RN(
        n2450), .Q(n477), .QN(n1980) );
  SDFFR_X2 shifted_reg_0_ ( .D(n1190), .SI(n1951), .SE(test_se), .CK(i_clk), 
        .RN(n2467), .Q(n2960), .QN(n3116) );
  SDFFR_X2 state_reg_reg_0_ ( .D(n1293), .SI(n2022), .SE(test_se), .CK(i_clk), 
        .RN(i_rst), .Q(n1954), .QN(n110) );
  SDFFR_X2 PR_reg_0_ ( .D(n52), .SI(n870), .SE(test_se), .CK(i_clk), .RN(n2459), .Q(n3053), .QN(n3025) );
  SDFFR_X2 ready_reg ( .D(n1230), .SI(n182), .SE(test_se), .CK(i_clk), .RN(
        n2462), .Q(ready), .QN(n171) );
  SDFFR_X2 reg_carry_reg ( .D(n1043), .SI(n2961), .SE(test_se), .CK(i_clk), 
        .RN(n2445), .Q(reg_carry), .QN(n395) );
  SDFFR_X2 DD_sign_reg ( .D(n1227), .SI(test_si1), .SE(test_se), .CK(i_clk), 
        .RN(n2445), .Q(n1955), .QN(n108) );
  SDFFR_X2 ct_1_en_1_reg ( .D(n1864), .SI(n3185), .SE(test_se), .CK(i_clk), 
        .RN(n2462), .Q(n3001), .QN(n169) );
  SDFFR_X2 ct_1_en_reg ( .D(n1113), .SI(n3001), .SE(test_se), .CK(i_clk), .RN(
        n2463), .Q(n1976), .QN(n109) );
  SDFFR_X2 shifted_1_reg_3_ ( .D(n2786), .SI(n1952), .SE(test_se), .CK(i_clk), 
        .RN(n2462), .Q(n1951), .QN(n172) );
  SDFFR_X2 shifted_1_reg_2_ ( .D(n2785), .SI(n1953), .SE(test_se), .CK(i_clk), 
        .RN(n2462), .Q(n1952), .QN(n173) );
  SDFFR_X2 shifted_1_reg_1_ ( .D(n2784), .SI(n1950), .SE(test_se), .CK(i_clk), 
        .RN(n2462), .Q(n1953), .QN(n174) );
  SDFFR_X2 shifted_1_reg_0_ ( .D(n2783), .SI(n2334), .SE(test_se), .CK(i_clk), 
        .RN(n2462), .Q(n1950), .QN(n175) );
  SDFFR_X2 DR_reg_30_ ( .D(n1125), .SI(n3182), .SE(test_se), .CK(i_clk), .RN(
        n2458), .Q(n3184), .QN(n121) );
  SDFFR_X2 DR_reg_29_ ( .D(n1126), .SI(n3180), .SE(test_se), .CK(i_clk), .RN(
        n2458), .Q(n3182), .QN(n122) );
  SDFFR_X2 DR_reg_28_ ( .D(n1127), .SI(n3178), .SE(test_se), .CK(i_clk), .RN(
        n2458), .Q(n3180), .QN(n123) );
  SDFFR_X2 DR_reg_27_ ( .D(n1128), .SI(n3176), .SE(test_se), .CK(i_clk), .RN(
        n2458), .Q(n3178), .QN(n124) );
  SDFFR_X2 DR_reg_26_ ( .D(n1129), .SI(n3174), .SE(test_se), .CK(i_clk), .RN(
        n2458), .Q(n3176), .QN(n125) );
  SDFFR_X2 DR_reg_25_ ( .D(n1130), .SI(n3172), .SE(test_se), .CK(i_clk), .RN(
        n2458), .Q(n3174), .QN(n126) );
  SDFFR_X2 DR_reg_24_ ( .D(n1131), .SI(n3170), .SE(test_se), .CK(i_clk), .RN(
        n2458), .Q(n3172), .QN(n127) );
  SDFFR_X2 DR_reg_23_ ( .D(n1132), .SI(n3168), .SE(test_se), .CK(i_clk), .RN(
        n2458), .Q(n3170), .QN(n128) );
  SDFFR_X2 DR_reg_22_ ( .D(n1133), .SI(n3166), .SE(test_se), .CK(i_clk), .RN(
        n2458), .Q(n3168), .QN(n129) );
  SDFFR_X2 DR_reg_10_ ( .D(n1145), .SI(n3142), .SE(test_se), .CK(i_clk), .RN(
        n2459), .Q(n3144), .QN(n141) );
  SDFFR_X2 DR_reg_31_ ( .D(n1124), .SI(n3184), .SE(test_se), .CK(i_clk), .RN(
        n2458), .Q(n3193), .QN(n119) );
  SDFFR_X2 DR_reg_21_ ( .D(n1134), .SI(n3164), .SE(test_se), .CK(i_clk), .RN(
        n2458), .Q(n3166), .QN(n130) );
  SDFFR_X2 DR_reg_20_ ( .D(n1135), .SI(n3162), .SE(test_se), .CK(i_clk), .RN(
        n2459), .Q(n3164), .QN(n131) );
  SDFFR_X2 DR_reg_19_ ( .D(n1136), .SI(n3160), .SE(test_se), .CK(i_clk), .RN(
        n2459), .Q(n3162), .QN(n132) );
  SDFFR_X2 DR_reg_18_ ( .D(n1137), .SI(n3158), .SE(test_se), .CK(i_clk), .RN(
        n2459), .Q(n3160), .QN(n133) );
  SDFFR_X2 DR_reg_17_ ( .D(n1138), .SI(n3156), .SE(test_se), .CK(i_clk), .RN(
        n2459), .Q(n3158), .QN(n134) );
  SDFFR_X2 DR_reg_16_ ( .D(n1139), .SI(n3154), .SE(test_se), .CK(i_clk), .RN(
        n2459), .Q(n3156), .QN(n135) );
  SDFFR_X2 DR_reg_15_ ( .D(n1140), .SI(n3152), .SE(test_se), .CK(i_clk), .RN(
        n2459), .Q(n3154), .QN(n136) );
  SDFFR_X2 DR_reg_14_ ( .D(n1141), .SI(n3150), .SE(test_se), .CK(i_clk), .RN(
        n2459), .Q(n3152), .QN(n137) );
  SDFFR_X2 DR_reg_13_ ( .D(n1142), .SI(n3148), .SE(test_se), .CK(i_clk), .RN(
        n2459), .Q(n3150), .QN(n138) );
  SDFFR_X2 DR_reg_12_ ( .D(n1143), .SI(n3146), .SE(test_se), .CK(i_clk), .RN(
        n2459), .Q(n3148), .QN(n139) );
  SDFFR_X2 DR_reg_11_ ( .D(n1144), .SI(n3144), .SE(test_se), .CK(i_clk), .RN(
        n2459), .Q(n3146), .QN(n140) );
  SDFFR_X2 DR_reg_9_ ( .D(n1146), .SI(n3140), .SE(test_se), .CK(i_clk), .RN(
        n2459), .Q(n3142), .QN(n142) );
  SDFFR_X2 DR_reg_8_ ( .D(n1147), .SI(n3138), .SE(test_se), .CK(i_clk), .RN(
        n2459), .Q(n3140), .QN(n143) );
  SDFFR_X2 DR_reg_7_ ( .D(n1148), .SI(n3136), .SE(test_se), .CK(i_clk), .RN(
        n2457), .Q(n3138), .QN(n111) );
  SDFFR_X2 DR_reg_6_ ( .D(n1149), .SI(n3134), .SE(test_se), .CK(i_clk), .RN(
        n2457), .Q(n3136), .QN(n112) );
  SDFFR_X2 DR_reg_5_ ( .D(n1150), .SI(n3131), .SE(test_se), .CK(i_clk), .RN(
        n2457), .Q(n3134), .QN(n113) );
  SDFFR_X2 DR_reg_4_ ( .D(n1151), .SI(n3128), .SE(test_se), .CK(i_clk), .RN(
        n2457), .Q(n3131), .QN(n114) );
  SDFFR_X2 DR_reg_3_ ( .D(n1152), .SI(n3125), .SE(test_se), .CK(i_clk), .RN(
        n2457), .Q(n3128), .QN(n115) );
  SDFFR_X2 DR_reg_2_ ( .D(n1153), .SI(n3122), .SE(test_se), .CK(i_clk), .RN(
        n2458), .Q(n3125), .QN(n116) );
  SDFFR_X2 DR_reg_1_ ( .D(n1154), .SI(n3187), .SE(test_se), .CK(i_clk), .RN(
        n2458), .Q(n3122), .QN(n117) );
  SDFFR_X2 DR_reg_0_ ( .D(n1155), .SI(n108), .SE(test_se), .CK(i_clk), .RN(
        n2458), .Q(n3187), .QN(n118) );
  SDFFR_X2 state_reg_reg_1_ ( .D(n2470), .SI(n1954), .SE(test_se), .CK(i_clk), 
        .RN(n2457), .Q(state_reg_1_0), .QN(test_so3) );
  SDFFR_X2 reg_b_reg_31_ ( .D(n4), .SI(reg_b[30]), .SE(test_se), .CK(i_clk), 
        .RN(n2447), .Q(reg_b[31]), .QN(n2961) );
  SDFFR_X2 nq_reg_30_ ( .D(n1075), .SI(nq[29]), .SE(test_se), .CK(i_clk), .RN(
        n2463), .Q(nq[30]), .QN(n183) );
  SDFFR_X2 nq_reg_29_ ( .D(n1076), .SI(n185), .SE(test_se), .CK(i_clk), .RN(
        n2463), .Q(nq[29]), .QN(n184) );
  SDFFR_X2 nq_reg_28_ ( .D(n1077), .SI(n186), .SE(test_se), .CK(i_clk), .RN(
        n2463), .Q(nq[28]), .QN(n185) );
  SDFFR_X2 nq_reg_27_ ( .D(n1078), .SI(n187), .SE(test_se), .CK(i_clk), .RN(
        n2463), .Q(nq[27]), .QN(n186) );
  SDFFR_X2 nq_reg_26_ ( .D(n1079), .SI(n188), .SE(test_se), .CK(i_clk), .RN(
        n2463), .Q(nq[26]), .QN(n187) );
  SDFFR_X2 nq_reg_25_ ( .D(n1080), .SI(n189), .SE(test_se), .CK(i_clk), .RN(
        n2463), .Q(nq[25]), .QN(n188) );
  SDFFR_X2 nq_reg_24_ ( .D(n1081), .SI(n220), .SE(test_se), .CK(i_clk), .RN(
        n2463), .Q(nq[24]), .QN(n189) );
  SDFFR_X2 nq_reg_7_ ( .D(n1098), .SI(n213), .SE(test_se), .CK(i_clk), .RN(
        n2465), .Q(nq[7]), .QN(n219) );
  SDFFR_X2 nq_reg_6_ ( .D(n1099), .SI(test_si2), .SE(test_se), .CK(i_clk), 
        .RN(n2465), .Q(nq[6]), .QN(n213) );
  SDFFR_X2 nq_reg_5_ ( .D(n1100), .SI(n2996), .SE(test_se), .CK(i_clk), .RN(
        n2465), .Q(nq[5]), .QN(n214) );
  SDFFR_X2 nq_reg_4_ ( .D(n1101), .SI(n2997), .SE(test_se), .CK(i_clk), .RN(
        n2465), .Q(n2996), .QN(n215) );
  SDFFR_X2 nq_reg_3_ ( .D(n1102), .SI(n2998), .SE(test_se), .CK(i_clk), .RN(
        n2465), .Q(n2997), .QN(n216) );
  SDFFR_X2 nq_reg_2_ ( .D(n1103), .SI(n2999), .SE(test_se), .CK(i_clk), .RN(
        n2465), .Q(n2998), .QN(n218) );
  SDFFR_X2 q_reg_30_ ( .D(n1044), .SI(q[29]), .SE(test_se), .CK(i_clk), .RN(
        n2463), .Q(q[30]), .QN(n182) );
  SDFFR_X2 nq_reg_8_ ( .D(n1097), .SI(n219), .SE(test_se), .CK(i_clk), .RN(
        n2466), .Q(nq[8]), .QN(n235) );
  SDFFR_X2 nq_reg_23_ ( .D(n1082), .SI(n221), .SE(test_se), .CK(i_clk), .RN(
        n2465), .Q(nq[23]), .QN(n220) );
  SDFFR_X2 nq_reg_22_ ( .D(n1083), .SI(n222), .SE(test_se), .CK(i_clk), .RN(
        n2465), .Q(nq[22]), .QN(n221) );
  SDFFR_X2 nq_reg_21_ ( .D(n1084), .SI(n223), .SE(test_se), .CK(i_clk), .RN(
        n2465), .Q(nq[21]), .QN(n222) );
  SDFFR_X2 nq_reg_20_ ( .D(n1085), .SI(n224), .SE(test_se), .CK(i_clk), .RN(
        n2465), .Q(nq[20]), .QN(n223) );
  SDFFR_X2 nq_reg_19_ ( .D(n1086), .SI(n225), .SE(test_se), .CK(i_clk), .RN(
        n2466), .Q(nq[19]), .QN(n224) );
  SDFFR_X2 nq_reg_18_ ( .D(n1087), .SI(n226), .SE(test_se), .CK(i_clk), .RN(
        n2466), .Q(nq[18]), .QN(n225) );
  SDFFR_X2 nq_reg_17_ ( .D(n1088), .SI(n227), .SE(test_se), .CK(i_clk), .RN(
        n2466), .Q(nq[17]), .QN(n226) );
  SDFFR_X2 nq_reg_16_ ( .D(n1089), .SI(n228), .SE(test_se), .CK(i_clk), .RN(
        n2466), .Q(nq[16]), .QN(n227) );
  SDFFR_X2 nq_reg_15_ ( .D(n1090), .SI(n229), .SE(test_se), .CK(i_clk), .RN(
        n2466), .Q(nq[15]), .QN(n228) );
  SDFFR_X2 nq_reg_14_ ( .D(n1091), .SI(n230), .SE(test_se), .CK(i_clk), .RN(
        n2466), .Q(nq[14]), .QN(n229) );
  SDFFR_X2 nq_reg_13_ ( .D(n1092), .SI(n231), .SE(test_se), .CK(i_clk), .RN(
        n2466), .Q(nq[13]), .QN(n230) );
  SDFFR_X2 nq_reg_12_ ( .D(n1093), .SI(n232), .SE(test_se), .CK(i_clk), .RN(
        n2466), .Q(nq[12]), .QN(n231) );
  SDFFR_X2 nq_reg_11_ ( .D(n1094), .SI(n233), .SE(test_se), .CK(i_clk), .RN(
        n2466), .Q(nq[11]), .QN(n232) );
  SDFFR_X2 nq_reg_10_ ( .D(n1095), .SI(n234), .SE(test_se), .CK(i_clk), .RN(
        n2466), .Q(nq[10]), .QN(n233) );
  SDFFR_X2 nq_reg_9_ ( .D(n1096), .SI(n235), .SE(test_se), .CK(i_clk), .RN(
        n2466), .Q(nq[9]), .QN(n234) );
  SDFFR_X2 q_reg_29_ ( .D(n1045), .SI(q[28]), .SE(test_se), .CK(i_clk), .RN(
        n2462), .Q(q[29]), .QN(n176) );
  SDFFR_X2 q_reg_28_ ( .D(n1046), .SI(test_si3), .SE(test_se), .CK(i_clk), 
        .RN(n2462), .Q(q[28]), .QN(n177) );
  SDFFR_X2 q_reg_27_ ( .D(n1047), .SI(q[26]), .SE(test_se), .CK(i_clk), .RN(
        n2462), .Q(q[27]), .QN(n178) );
  SDFFR_X2 q_reg_26_ ( .D(n1048), .SI(q[25]), .SE(test_se), .CK(i_clk), .RN(
        n2462), .Q(q[26]), .QN(n179) );
  SDFFR_X2 q_reg_25_ ( .D(n1049), .SI(q[24]), .SE(test_se), .CK(i_clk), .RN(
        n2462), .Q(q[25]), .QN(n180) );
  SDFFR_X2 q_reg_24_ ( .D(n1050), .SI(q[23]), .SE(test_se), .CK(i_clk), .RN(
        n2462), .Q(q[24]), .QN(n181) );
  SDFFR_X2 q_reg_1_ ( .D(n1073), .SI(n398), .SE(test_se), .CK(i_clk), .RN(
        n2464), .Q(q[1]), .QN(n195) );
  SDFFR_X2 q_reg_0_ ( .D(n1074), .SI(o_remainder[30]), .SE(test_se), .CK(i_clk), .RN(n2446), .Q(q[0]), .QN(n398) );
  SDFFR_X2 q_reg_7_ ( .D(n1067), .SI(q[6]), .SE(test_se), .CK(i_clk), .RN(
        n2463), .Q(q[7]), .QN(n190) );
  SDFFR_X2 q_reg_6_ ( .D(n1068), .SI(q[5]), .SE(test_se), .CK(i_clk), .RN(
        n2463), .Q(q[6]), .QN(n191) );
  SDFFR_X2 q_reg_5_ ( .D(n1069), .SI(q[4]), .SE(test_se), .CK(i_clk), .RN(
        n2464), .Q(q[5]), .QN(n196) );
  SDFFR_X2 q_reg_4_ ( .D(n1070), .SI(q[3]), .SE(test_se), .CK(i_clk), .RN(
        n2463), .Q(q[4]), .QN(n192) );
  SDFFR_X2 q_reg_3_ ( .D(n1071), .SI(n194), .SE(test_se), .CK(i_clk), .RN(
        n2463), .Q(q[3]), .QN(n193) );
  SDFFR_X2 q_reg_2_ ( .D(n1072), .SI(n195), .SE(test_se), .CK(i_clk), .RN(
        n2463), .Q(q[2]), .QN(n194) );
  SDFFR_X2 q_reg_23_ ( .D(n1051), .SI(q[22]), .SE(test_se), .CK(i_clk), .RN(
        n2464), .Q(q[23]), .QN(n201) );
  SDFFR_X2 q_reg_22_ ( .D(n1052), .SI(q[21]), .SE(test_se), .CK(i_clk), .RN(
        n2464), .Q(q[22]), .QN(n202) );
  SDFFR_X2 q_reg_21_ ( .D(n1053), .SI(q[20]), .SE(test_se), .CK(i_clk), .RN(
        n2464), .Q(q[21]), .QN(n203) );
  SDFFR_X2 q_reg_20_ ( .D(n1054), .SI(q[19]), .SE(test_se), .CK(i_clk), .RN(
        n2464), .Q(q[20]), .QN(n204) );
  SDFFR_X2 q_reg_19_ ( .D(n1055), .SI(q[18]), .SE(test_se), .CK(i_clk), .RN(
        n2464), .Q(q[19]), .QN(n205) );
  SDFFR_X2 q_reg_18_ ( .D(n1056), .SI(q[17]), .SE(test_se), .CK(i_clk), .RN(
        n2464), .Q(q[18]), .QN(n206) );
  SDFFR_X2 q_reg_17_ ( .D(n1057), .SI(q[16]), .SE(test_se), .CK(i_clk), .RN(
        n2464), .Q(q[17]), .QN(n207) );
  SDFFR_X2 q_reg_16_ ( .D(n1058), .SI(q[15]), .SE(test_se), .CK(i_clk), .RN(
        n2464), .Q(q[16]), .QN(n208) );
  SDFFR_X2 q_reg_15_ ( .D(n1059), .SI(q[14]), .SE(test_se), .CK(i_clk), .RN(
        n2465), .Q(q[15]), .QN(n209) );
  SDFFR_X2 q_reg_14_ ( .D(n1060), .SI(q[13]), .SE(test_se), .CK(i_clk), .RN(
        n2465), .Q(q[14]), .QN(n210) );
  SDFFR_X2 q_reg_13_ ( .D(n1061), .SI(q[12]), .SE(test_se), .CK(i_clk), .RN(
        n2465), .Q(q[13]), .QN(n211) );
  SDFFR_X2 q_reg_12_ ( .D(n1062), .SI(q[11]), .SE(test_se), .CK(i_clk), .RN(
        n2465), .Q(q[12]), .QN(n212) );
  SDFFR_X2 q_reg_11_ ( .D(n1063), .SI(q[10]), .SE(test_se), .CK(i_clk), .RN(
        n2464), .Q(q[11]), .QN(n197) );
  SDFFR_X2 q_reg_10_ ( .D(n1064), .SI(q[9]), .SE(test_se), .CK(i_clk), .RN(
        n2464), .Q(q[10]), .QN(n198) );
  SDFFR_X2 q_reg_9_ ( .D(n1065), .SI(q[8]), .SE(test_se), .CK(i_clk), .RN(
        n2464), .Q(q[9]), .QN(n199) );
  SDFFR_X2 q_reg_8_ ( .D(n1066), .SI(q[7]), .SE(test_se), .CK(i_clk), .RN(
        n2464), .Q(q[8]), .QN(n200) );
  SDFFR_X2 reg_b_reg_0_ ( .D(n1292), .SI(n2968), .SE(test_se), .CK(i_clk), 
        .RN(n2467), .Q(reg_b[0]), .QN(n281) );
  SDFFR_X2 reg_a_reg_0_ ( .D(n1042), .SI(ready), .SE(test_se), .CK(i_clk), 
        .RN(n2453), .Q(reg_a[0]), .QN(n2993) );
  SDFFR_X2 reg_a_reg_1_ ( .D(n1041), .SI(n2993), .SE(test_se), .CK(i_clk), 
        .RN(n2453), .Q(reg_a[1]), .QN(n2992) );
  SDFFR_X2 reg_a_reg_3_ ( .D(n1039), .SI(n492), .SE(test_se), .CK(i_clk), .RN(
        n2453), .Q(reg_a[3]), .QN(n2991) );
  SDFFR_X2 state_reg_5_ ( .D(n1229), .SI(state[4]), .SE(test_se), .CK(i_clk), 
        .RN(n2466), .Q(n2022), .QN(n2335) );
  SDFFR_X2 state_reg_4_ ( .D(n1192), .SI(n241), .SE(test_se), .CK(i_clk), .RN(
        n2467), .Q(state[4]), .QN(n240) );
  SDFFR_X2 state_reg_3_ ( .D(n1225), .SI(n238), .SE(test_se), .CK(i_clk), .RN(
        n2467), .Q(state[3]), .QN(n241) );
  SDFFR_X2 state_reg_2_ ( .D(n1226), .SI(n239), .SE(test_se), .CK(i_clk), .RN(
        n2466), .Q(state[2]), .QN(n238) );
  SDFFR_X2 state_reg_1_ ( .D(n1228), .SI(n105), .SE(test_se), .CK(i_clk), .RN(
        n2467), .Q(state[1]), .QN(n239) );
  SDFFR_X2 reg_b_reg_5_ ( .D(n1287), .SI(n274), .SE(test_se), .CK(i_clk), .RN(
        n2467), .Q(reg_b[5]), .QN(n2965) );
  SDFFR_X2 reg_b_reg_1_ ( .D(n1291), .SI(n281), .SE(test_se), .CK(i_clk), .RN(
        n2467), .Q(reg_b[1]), .QN(n2967) );
  SDFFR_X2 sdata_reg_0_ ( .D(n1186), .SI(n395), .SE(test_se), .CK(i_clk), .RN(
        n2468), .Q(sdata[0]), .QN(n298) );
  SDFFR_X2 reg_b_reg_3_ ( .D(n1289), .SI(reg_b[2]), .SE(test_se), .CK(i_clk), 
        .RN(n2467), .Q(reg_b[3]), .QN(n2966) );
  SDFFR_X2 reg_a_reg_2_ ( .D(n1040), .SI(n2992), .SE(test_se), .CK(i_clk), 
        .RN(n2453), .Q(reg_a[2]), .QN(n492) );
  SDFFR_X2 reg_b_reg_11_ ( .D(n1281), .SI(n488), .SE(test_se), .CK(i_clk), 
        .RN(n2450), .Q(reg_b[11]), .QN(n480) );
  SDFFR_X2 reg_b_reg_9_ ( .D(n1283), .SI(n484), .SE(test_se), .CK(i_clk), .RN(
        n2451), .Q(reg_b[9]), .QN(n483) );
  SDFFR_X2 reg_b_reg_7_ ( .D(n1285), .SI(n2964), .SE(test_se), .CK(i_clk), 
        .RN(n2451), .Q(reg_b[7]), .QN(n486) );
  SDFFR_X2 reg_a_reg_31_ ( .D(n1011), .SI(n2969), .SE(test_se), .CK(i_clk), 
        .RN(n2452), .Q(reg_a[31]), .QN(n2968) );
  SDFFR_X2 reg_a_reg_6_ ( .D(n1036), .SI(n2990), .SE(test_se), .CK(i_clk), 
        .RN(n2454), .Q(reg_a[6]), .QN(n497) );
  SDFFR_X2 reg_a_reg_4_ ( .D(n1038), .SI(n2991), .SE(test_se), .CK(i_clk), 
        .RN(n2453), .Q(reg_a[4]), .QN(n491) );
  SDFFR_X2 reg_a_reg_12_ ( .D(n1030), .SI(n2985), .SE(test_se), .CK(i_clk), 
        .RN(n2454), .Q(reg_a[12]), .QN(n2984) );
  SDFFR_X2 reg_a_reg_10_ ( .D(n1032), .SI(n2987), .SE(test_se), .CK(i_clk), 
        .RN(n2454), .Q(reg_a[10]), .QN(n2986) );
  SDFFR_X2 reg_a_reg_8_ ( .D(n1034), .SI(n2989), .SE(test_se), .CK(i_clk), 
        .RN(n2454), .Q(reg_a[8]), .QN(n2988) );
  SDFFR_X2 reg_a_reg_7_ ( .D(n1035), .SI(n497), .SE(test_se), .CK(i_clk), .RN(
        n2454), .Q(reg_a[7]), .QN(n2989) );
  SDFFR_X2 reg_a_reg_5_ ( .D(n1037), .SI(reg_a[4]), .SE(test_se), .CK(i_clk), 
        .RN(n2454), .Q(reg_a[5]), .QN(n2990) );
  SDFFR_X2 reg_a_reg_13_ ( .D(n1029), .SI(n2984), .SE(test_se), .CK(i_clk), 
        .RN(n2454), .Q(reg_a[13]), .QN(n2983) );
  SDFFR_X2 reg_a_reg_11_ ( .D(n1031), .SI(n2986), .SE(test_se), .CK(i_clk), 
        .RN(n2454), .Q(reg_a[11]), .QN(n2985) );
  SDFFR_X2 reg_a_reg_9_ ( .D(n1033), .SI(n2988), .SE(test_se), .CK(i_clk), 
        .RN(n2454), .Q(reg_a[9]), .QN(n2987) );
  SDFFR_X2 reg_b_reg_4_ ( .D(n1288), .SI(n2966), .SE(test_se), .CK(i_clk), 
        .RN(n2467), .Q(reg_b[4]), .QN(n274) );
  SDFFR_X2 reg_b_reg_2_ ( .D(n1290), .SI(n2967), .SE(test_se), .CK(i_clk), 
        .RN(n2467), .Q(reg_b[2]), .QN(n279) );
  SDFFR_X2 PR_reg_2_ ( .D(n56), .SI(n3024), .SE(test_se), .CK(i_clk), .RN(
        n2462), .Q(n3123), .QN(n3023) );
  SDFFR_X2 PR_reg_1_ ( .D(n51), .SI(n3025), .SE(test_se), .CK(i_clk), .RN(
        n2461), .Q(n3120), .QN(n3024) );
  SDFFR_X2 reg_b_reg_13_ ( .D(n1279), .SI(n489), .SE(test_se), .CK(i_clk), 
        .RN(n2454), .Q(reg_b[13]), .QN(n493) );
  SDFFR_X2 reg_b_reg_12_ ( .D(n1280), .SI(n480), .SE(test_se), .CK(i_clk), 
        .RN(n2452), .Q(reg_b[12]), .QN(n489) );
  SDFFR_X2 reg_b_reg_10_ ( .D(n1282), .SI(n483), .SE(test_se), .CK(i_clk), 
        .RN(n2452), .Q(reg_b[10]), .QN(n488) );
  SDFFR_X2 reg_b_reg_8_ ( .D(n1284), .SI(n486), .SE(test_se), .CK(i_clk), .RN(
        n2451), .Q(reg_b[8]), .QN(n484) );
  SDFFR_X2 reg_b_reg_6_ ( .D(n1286), .SI(n2965), .SE(test_se), .CK(i_clk), 
        .RN(n2451), .Q(n2964), .QN(n487) );
  SDFFR_X2 reg_a_reg_15_ ( .D(n1027), .SI(n500), .SE(test_se), .CK(i_clk), 
        .RN(n2455), .Q(reg_a[15]), .QN(n2982) );
  SDFFR_X2 reg_a_reg_14_ ( .D(n1028), .SI(n2983), .SE(test_se), .CK(i_clk), 
        .RN(n2454), .Q(reg_a[14]), .QN(n500) );
  SDFFR_X2 reg_b_reg_14_ ( .D(n1278), .SI(n493), .SE(test_se), .CK(i_clk), 
        .RN(n2454), .Q(reg_b[14]), .QN(n499) );
  SDFFR_X2 sdata_reg_31_ ( .D(n1296), .SI(sdata[30]), .SE(test_se), .CK(i_clk), 
        .RN(n2457), .Q(n2019), .QN(n2334) );
  SDFFR_X2 reg_a_reg_17_ ( .D(n1025), .SI(n2981), .SE(test_se), .CK(i_clk), 
        .RN(n2455), .Q(reg_a[17]), .QN(n2980) );
  SDFFR_X2 reg_a_reg_16_ ( .D(n1026), .SI(n2982), .SE(test_se), .CK(i_clk), 
        .RN(n2455), .Q(reg_a[16]), .QN(n2981) );
  SDFFR_X2 reg_b_reg_15_ ( .D(n1277), .SI(n499), .SE(test_se), .CK(i_clk), 
        .RN(n2455), .Q(reg_b[15]), .QN(n502) );
  SDFFR_X2 sdata_reg_2_ ( .D(n1184), .SI(n345), .SE(test_se), .CK(i_clk), .RN(
        n2469), .Q(sdata[2]), .QN(n390) );
  SDFFR_X2 sdata_reg_1_ ( .D(n1185), .SI(n298), .SE(test_se), .CK(i_clk), .RN(
        n2468), .Q(sdata[1]), .QN(n345) );
  SDFFR_X2 reg_b_reg_16_ ( .D(n1276), .SI(reg_b[15]), .SE(test_se), .CK(i_clk), 
        .RN(n2455), .Q(reg_b[16]), .QN(n505) );
  SDFFR_X2 PR_reg_3_ ( .D(n55), .SI(n3023), .SE(test_se), .CK(i_clk), .RN(
        n2462), .Q(n3126), .QN(n3022) );
  SDFFR_X2 PR_reg_4_ ( .D(n54), .SI(n3022), .SE(test_se), .CK(i_clk), .RN(
        n2461), .Q(n3129), .QN(n3021) );
  SDFFR_X2 reg_a_reg_19_ ( .D(n1023), .SI(n2979), .SE(test_se), .CK(i_clk), 
        .RN(n2455), .Q(reg_a[19]), .QN(n2978) );
  SDFFR_X2 reg_a_reg_18_ ( .D(n1024), .SI(n2980), .SE(test_se), .CK(i_clk), 
        .RN(n2455), .Q(reg_a[18]), .QN(n2979) );
  SDFFR_X2 reg_b_reg_17_ ( .D(n1275), .SI(n505), .SE(test_se), .CK(i_clk), 
        .RN(n2455), .Q(reg_b[17]), .QN(n510) );
  SDFFR_X2 reg_b_reg_18_ ( .D(n1274), .SI(n510), .SE(test_se), .CK(i_clk), 
        .RN(n2455), .Q(reg_b[18]), .QN(n513) );
  SDFFR_X2 sdata_reg_3_ ( .D(n1183), .SI(n390), .SE(test_se), .CK(i_clk), .RN(
        n2469), .Q(sdata[3]), .QN(n387) );
  SDFFR_X2 reg_a_reg_21_ ( .D(n1021), .SI(n2977), .SE(test_se), .CK(i_clk), 
        .RN(n2456), .Q(reg_a[21]), .QN(n2976) );
  SDFFR_X2 sdata_reg_4_ ( .D(n1182), .SI(n387), .SE(test_se), .CK(i_clk), .RN(
        n2469), .Q(sdata[4]), .QN(n386) );
  SDFFR_X2 reg_a_reg_20_ ( .D(n1022), .SI(n2978), .SE(test_se), .CK(i_clk), 
        .RN(n2455), .Q(reg_a[20]), .QN(n2977) );
  SDFFR_X2 reg_b_reg_19_ ( .D(n1273), .SI(n513), .SE(test_se), .CK(i_clk), 
        .RN(n2455), .Q(reg_b[19]), .QN(n511) );
  SDFFR_X2 reg_b_reg_20_ ( .D(n1272), .SI(n511), .SE(test_se), .CK(i_clk), 
        .RN(n2455), .Q(reg_b[20]), .QN(n514) );
  SDFFR_X2 reg_a_reg_23_ ( .D(n1019), .SI(n2975), .SE(test_se), .CK(i_clk), 
        .RN(n2456), .Q(reg_a[23]), .QN(n2974) );
  SDFFR_X2 reg_a_reg_22_ ( .D(n1020), .SI(n2976), .SE(test_se), .CK(i_clk), 
        .RN(n2456), .Q(reg_a[22]), .QN(n2975) );
  SDFFR_X2 PR_reg_30_ ( .D(n838), .SI(n3002), .SE(test_se), .CK(i_clk), .RN(
        n2460), .Q(n1977), .QN(n154) );
  SDFFR_X2 reg_b_reg_21_ ( .D(n1271), .SI(n514), .SE(test_se), .CK(i_clk), 
        .RN(n2455), .Q(reg_b[21]), .QN(n517) );
  SDFFR_X2 PR_reg_6_ ( .D(n862), .SI(n3020), .SE(test_se), .CK(i_clk), .RN(
        n2461), .Q(n3019), .QN(n165) );
  SDFFR_X2 PR_reg_7_ ( .D(n861), .SI(n3019), .SE(test_se), .CK(i_clk), .RN(
        n2461), .Q(n3018), .QN(n164) );
  SDFFR_X2 reg_b_reg_22_ ( .D(n1270), .SI(reg_b[21]), .SE(test_se), .CK(i_clk), 
        .RN(n2455), .Q(reg_b[22]), .QN(n518) );
  SDFFR_X2 PR_reg_5_ ( .D(n53), .SI(n3021), .SE(test_se), .CK(i_clk), .RN(
        n2461), .Q(n3132), .QN(n3020) );
  SDFFR_X2 reg_a_reg_24_ ( .D(n1018), .SI(n2974), .SE(test_se), .CK(i_clk), 
        .RN(n2456), .Q(reg_a[24]), .QN(n2973) );
  SDFFR_X2 PR_reg_24_ ( .D(n47), .SI(n3005), .SE(test_se), .CK(i_clk), .RN(
        n2461), .Q(n1957), .QN(n158) );
  SDFFR_X2 PR_reg_22_ ( .D(n48), .SI(n3006), .SE(test_se), .CK(i_clk), .RN(
        n2460), .Q(n1959), .QN(n153) );
  SDFFR_X2 PR_reg_20_ ( .D(n49), .SI(n3007), .SE(test_se), .CK(i_clk), .RN(
        n2461), .Q(n1947), .QN(n160) );
  SDFFR_X2 PR_reg_18_ ( .D(n50), .SI(n3008), .SE(test_se), .CK(i_clk), .RN(
        n2461), .Q(n1949), .QN(n163) );
  SDFFR_X2 PR_reg_28_ ( .D(n840), .SI(n1966), .SE(test_se), .CK(i_clk), .RN(
        n2461), .Q(n3003), .QN(n168) );
  SDFFR_X2 PR_reg_29_ ( .D(n839), .SI(n3003), .SE(test_se), .CK(i_clk), .RN(
        n2460), .Q(n3002), .QN(n155) );
  SDFFR_X2 reg_a_reg_26_ ( .D(n1016), .SI(n2972), .SE(test_se), .CK(i_clk), 
        .RN(n2456), .Q(reg_a[26]), .QN(n526) );
  SDFFR_X2 reg_a_reg_25_ ( .D(n1017), .SI(n2973), .SE(test_se), .CK(i_clk), 
        .RN(n2456), .Q(reg_a[25]), .QN(n2972) );
  SDFFR_X2 PR_reg_8_ ( .D(n860), .SI(n3018), .SE(test_se), .CK(i_clk), .RN(
        n2461), .Q(n3017), .QN(n166) );
  SDFFR_X2 PR_reg_14_ ( .D(n854), .SI(n3012), .SE(test_se), .CK(i_clk), .RN(
        n2460), .Q(n3011), .QN(n149) );
  SDFFR_X2 PR_reg_13_ ( .D(n855), .SI(n3013), .SE(test_se), .CK(i_clk), .RN(
        n2460), .Q(n3012), .QN(n145) );
  SDFFR_X2 PR_reg_12_ ( .D(n856), .SI(n3014), .SE(test_se), .CK(i_clk), .RN(
        n2460), .Q(n3013), .QN(n146) );
  SDFFR_X2 PR_reg_11_ ( .D(n857), .SI(n3015), .SE(test_se), .CK(i_clk), .RN(
        n2460), .Q(n3014), .QN(n147) );
  SDFFR_X2 PR_reg_10_ ( .D(n858), .SI(n3016), .SE(test_se), .CK(i_clk), .RN(
        n2460), .Q(n3015), .QN(n150) );
  SDFFR_X2 PR_reg_9_ ( .D(n859), .SI(n3017), .SE(test_se), .CK(i_clk), .RN(
        n2461), .Q(n3016), .QN(n167) );
  SDFFR_X2 PR_reg_16_ ( .D(n852), .SI(n3010), .SE(test_se), .CK(i_clk), .RN(
        n2460), .Q(n3009), .QN(n148) );
  SDFFR_X2 PR_reg_17_ ( .D(n851), .SI(n3009), .SE(test_se), .CK(i_clk), .RN(
        n2461), .Q(n3008), .QN(n162) );
  SDFFR_X2 PR_reg_15_ ( .D(n853), .SI(n3011), .SE(test_se), .CK(i_clk), .RN(
        n2460), .Q(n3010), .QN(n144) );
  SDFFR_X2 PR_reg_26_ ( .D(n46), .SI(n3004), .SE(test_se), .CK(i_clk), .RN(
        n2460), .Q(n1967), .QN(n151) );
  SDFFR_X2 sdata_reg_30_ ( .D(n1156), .SI(sdata[29]), .SE(test_se), .CK(i_clk), 
        .RN(n2457), .Q(sdata[30]), .QN(n534) );
  SDFFR_X2 PR_reg_25_ ( .D(n843), .SI(n1957), .SE(test_se), .CK(i_clk), .RN(
        n2460), .Q(n3004), .QN(n157) );
  SDFFR_X2 PR_reg_23_ ( .D(n845), .SI(n1959), .SE(test_se), .CK(i_clk), .RN(
        n2460), .Q(n3005), .QN(n152) );
  SDFFR_X2 PR_reg_21_ ( .D(n847), .SI(n1947), .SE(test_se), .CK(i_clk), .RN(
        n2461), .Q(n3006), .QN(n159) );
  SDFFR_X2 PR_reg_19_ ( .D(n849), .SI(n1949), .SE(test_se), .CK(i_clk), .RN(
        n2461), .Q(n3007), .QN(n161) );
  SDFFR_X2 PR_reg_27_ ( .D(n45), .SI(n1967), .SE(test_se), .CK(i_clk), .RN(
        n2460), .Q(n1966), .QN(n156) );
  SDFFR_X2 reg_b_reg_23_ ( .D(n1269), .SI(n518), .SE(test_se), .CK(i_clk), 
        .RN(n2456), .Q(reg_b[23]), .QN(n519) );
  SDFFR_X2 sdata_reg_5_ ( .D(n1181), .SI(n386), .SE(test_se), .CK(i_clk), .RN(
        n2469), .Q(sdata[5]), .QN(n385) );
  SDFFR_X2 sdata_reg_6_ ( .D(n1180), .SI(n385), .SE(test_se), .CK(i_clk), .RN(
        n2469), .Q(sdata[6]), .QN(n388) );
  SDFFR_X2 reg_b_reg_24_ ( .D(n1268), .SI(n519), .SE(test_se), .CK(i_clk), 
        .RN(n2456), .Q(reg_b[24]), .QN(n522) );
  SDFFR_X2 sdata_reg_26_ ( .D(n1160), .SI(sdata[25]), .SE(test_se), .CK(i_clk), 
        .RN(n2468), .Q(sdata[26]), .QN(n372) );
  SDFFR_X2 sdata_reg_7_ ( .D(n1179), .SI(n388), .SE(test_se), .CK(i_clk), .RN(
        n2469), .Q(sdata[7]), .QN(n389) );
  SDFFR_X2 sdata_reg_22_ ( .D(n1164), .SI(n377), .SE(test_se), .CK(i_clk), 
        .RN(n2469), .Q(sdata[22]), .QN(n376) );
  SDFFR_X2 sdata_reg_20_ ( .D(n1166), .SI(n379), .SE(test_se), .CK(i_clk), 
        .RN(n2469), .Q(sdata[20]), .QN(n378) );
  SDFFR_X2 sdata_reg_18_ ( .D(n1168), .SI(n380), .SE(test_se), .CK(i_clk), 
        .RN(n2469), .Q(sdata[18]), .QN(n381) );
  SDFFR_X2 sdata_reg_23_ ( .D(n1163), .SI(sdata[22]), .SE(test_se), .CK(i_clk), 
        .RN(n2468), .Q(sdata[23]), .QN(n375) );
  SDFFR_X2 sdata_reg_21_ ( .D(n1165), .SI(n378), .SE(test_se), .CK(i_clk), 
        .RN(n2469), .Q(sdata[21]), .QN(n377) );
  SDFFR_X2 sdata_reg_19_ ( .D(n1167), .SI(n381), .SE(test_se), .CK(i_clk), 
        .RN(n2469), .Q(sdata[19]), .QN(n379) );
  SDFFR_X2 sdata_reg_24_ ( .D(n1162), .SI(sdata[23]), .SE(test_se), .CK(i_clk), 
        .RN(n2468), .Q(sdata[24]), .QN(n374) );
  SDFFR_X2 sdata_reg_25_ ( .D(n1161), .SI(sdata[24]), .SE(test_se), .CK(i_clk), 
        .RN(n2468), .Q(sdata[25]), .QN(n373) );
  SDFFR_X2 sdata_reg_10_ ( .D(n1176), .SI(n392), .SE(test_se), .CK(i_clk), 
        .RN(n2468), .Q(sdata[10]), .QN(n342) );
  SDFFR_X2 sdata_reg_9_ ( .D(n1177), .SI(n391), .SE(test_se), .CK(i_clk), .RN(
        i_rst), .Q(sdata[9]), .QN(n392) );
  SDFFR_X2 sdata_reg_8_ ( .D(n1178), .SI(n389), .SE(test_se), .CK(i_clk), .RN(
        n2469), .Q(sdata[8]), .QN(n391) );
  SDFFR_X2 sdata_reg_16_ ( .D(n1170), .SI(n336), .SE(test_se), .CK(i_clk), 
        .RN(n2468), .Q(sdata[16]), .QN(n335) );
  SDFFR_X2 sdata_reg_15_ ( .D(n1171), .SI(n337), .SE(test_se), .CK(i_clk), 
        .RN(n2468), .Q(sdata[15]), .QN(n336) );
  SDFFR_X2 sdata_reg_14_ ( .D(n1172), .SI(n338), .SE(test_se), .CK(i_clk), 
        .RN(n2468), .Q(sdata[14]), .QN(n337) );
  SDFFR_X2 sdata_reg_13_ ( .D(n1173), .SI(n339), .SE(test_se), .CK(i_clk), 
        .RN(n2468), .Q(sdata[13]), .QN(n338) );
  SDFFR_X2 sdata_reg_12_ ( .D(n1174), .SI(n322), .SE(test_se), .CK(i_clk), 
        .RN(n2468), .Q(sdata[12]), .QN(n339) );
  SDFFR_X2 sdata_reg_11_ ( .D(n1175), .SI(n342), .SE(test_se), .CK(i_clk), 
        .RN(n2468), .Q(sdata[11]), .QN(n322) );
  SDFFR_X2 sdata_reg_17_ ( .D(n1169), .SI(n335), .SE(test_se), .CK(i_clk), 
        .RN(n2469), .Q(sdata[17]), .QN(n380) );
  SDFFR_X2 sdata_reg_29_ ( .D(n1157), .SI(sdata[28]), .SE(test_se), .CK(i_clk), 
        .RN(n2469), .Q(sdata[29]), .QN(n384) );
  SDFFR_X2 sdata_reg_28_ ( .D(n1158), .SI(sdata[27]), .SE(test_se), .CK(i_clk), 
        .RN(n2457), .Q(sdata[28]), .QN(n535) );
  SDFFR_X2 sdata_reg_27_ ( .D(n1159), .SI(sdata[26]), .SE(test_se), .CK(i_clk), 
        .RN(n2468), .Q(sdata[27]), .QN(n370) );
  SDFFR_X2 reg_a_reg_27_ ( .D(n1015), .SI(n526), .SE(test_se), .CK(i_clk), 
        .RN(n2456), .Q(reg_a[27]), .QN(n2971) );
  SDFFR_X2 reg_a_reg_28_ ( .D(n1014), .SI(n2971), .SE(test_se), .CK(i_clk), 
        .RN(n2457), .Q(reg_a[28]), .QN(n536) );
  SDFFR_X2 reg_a_reg_29_ ( .D(n1013), .SI(n536), .SE(test_se), .CK(i_clk), 
        .RN(n2456), .Q(reg_a[29]), .QN(n2970) );
  SDFFR_X2 reg_b_reg_25_ ( .D(n1267), .SI(n522), .SE(test_se), .CK(i_clk), 
        .RN(n2456), .Q(reg_b[25]), .QN(n524) );
  SDFFR_X2 reg_b_reg_26_ ( .D(n1266), .SI(reg_b[25]), .SE(test_se), .CK(i_clk), 
        .RN(n2456), .Q(n2963), .QN(n525) );
  SDFFR_X2 reg_a_reg_30_ ( .D(n1012), .SI(n2970), .SE(test_se), .CK(i_clk), 
        .RN(n2456), .Q(reg_a[30]), .QN(n2969) );
  SDFFR_X2 reg_b_reg_27_ ( .D(n1265), .SI(n2963), .SE(test_se), .CK(i_clk), 
        .RN(n2456), .Q(reg_b[27]), .QN(n529) );
  SDFFR_X2 reg_b_reg_28_ ( .D(n1264), .SI(reg_b[27]), .SE(test_se), .CK(i_clk), 
        .RN(n2457), .Q(n2962), .QN(n531) );
  SDFFR_X2 reg_b_reg_29_ ( .D(n1263), .SI(n2962), .SE(test_se), .CK(i_clk), 
        .RN(n2457), .Q(reg_b[29]), .QN(n537) );
  SDFFR_X2 reg_b_reg_30_ ( .D(n1297), .SI(n537), .SE(test_se), .CK(i_clk), 
        .RN(n2457), .Q(reg_b[30]), .QN(n538) );
  AND2_X4 U1940 ( .A1(n949), .A2(n948), .ZN(n2016) );
  AND4_X4 U1941 ( .A1(n2394), .A2(n68), .A3(n754), .A4(n2428), .ZN(n2017) );
  AND2_X4 U1942 ( .A1(n948), .A2(n445), .ZN(n2018) );
  XOR2_X2 U1943 ( .A(n534), .B(n2019), .Z(n2020) );
  OR2_X4 U1944 ( .A1(n1551), .A2(n1552), .ZN(n2021) );
  NOR2_X2 U1945 ( .A1(n110), .A2(state_reg_1_0), .ZN(n2023) );
  OR2_X4 U1946 ( .A1(n1855), .A2(n719), .ZN(n2024) );
  OR2_X4 U1947 ( .A1(n1869), .A2(n719), .ZN(n2025) );
  AND2_X4 U1948 ( .A1(n37), .A2(n1816), .ZN(n2026) );
  INV_X4 U2236 ( .A(n2314), .ZN(n2381) );
  INV_X4 U2237 ( .A(n2314), .ZN(n2382) );
  INV_X4 U2238 ( .A(n2443), .ZN(n2442) );
  AND2_X2 U2239 ( .A1(n1301), .A2(n2440), .ZN(n2314) );
  INV_X4 U2240 ( .A(n2315), .ZN(n2376) );
  INV_X4 U2241 ( .A(n2315), .ZN(n2375) );
  INV_X4 U2242 ( .A(n2315), .ZN(n2377) );
  INV_X4 U2243 ( .A(n2322), .ZN(n2443) );
  INV_X4 U2244 ( .A(n2444), .ZN(n2441) );
  INV_X4 U2245 ( .A(n2322), .ZN(n2444) );
  INV_X4 U2246 ( .A(n2390), .ZN(n2388) );
  INV_X4 U2247 ( .A(n2390), .ZN(n2389) );
  INV_X4 U2248 ( .A(n1318), .ZN(n361) );
  OR2_X2 U2249 ( .A1(n2387), .A2(n2438), .ZN(n2315) );
  INV_X4 U2250 ( .A(n2316), .ZN(n2373) );
  INV_X4 U2251 ( .A(n2317), .ZN(n2370) );
  INV_X4 U2252 ( .A(n2317), .ZN(n2371) );
  INV_X4 U2253 ( .A(n2316), .ZN(n2374) );
  INV_X4 U2254 ( .A(n1575), .ZN(n2440) );
  INV_X4 U2255 ( .A(n1575), .ZN(n2439) );
  INV_X4 U2256 ( .A(n2380), .ZN(n2378) );
  INV_X4 U2257 ( .A(n2380), .ZN(n2379) );
  INV_X4 U2258 ( .A(n2317), .ZN(n2372) );
  INV_X4 U2259 ( .A(n634), .ZN(n42) );
  INV_X4 U2260 ( .A(n2361), .ZN(n2362) );
  INV_X4 U2261 ( .A(n966), .ZN(n2390) );
  INV_X4 U2262 ( .A(n966), .ZN(n2391) );
  NAND2_X2 U2263 ( .A1(n364), .A2(n1551), .ZN(n1318) );
  AND2_X2 U2264 ( .A1(n2372), .A2(n2384), .ZN(n2316) );
  NAND3_X2 U2265 ( .A1(n1318), .A2(n2021), .A3(n1319), .ZN(n723) );
  AND2_X2 U2266 ( .A1(n367), .A2(n2439), .ZN(n2317) );
  NAND3_X2 U2267 ( .A1(n501), .A2(n955), .A3(n951), .ZN(n943) );
  INV_X4 U2268 ( .A(n1301), .ZN(n2380) );
  INV_X4 U2269 ( .A(n2021), .ZN(n2343) );
  INV_X4 U2270 ( .A(n978), .ZN(n2437) );
  INV_X4 U2271 ( .A(n2020), .ZN(n2386) );
  INV_X4 U2272 ( .A(n978), .ZN(n2436) );
  INV_X4 U2273 ( .A(n2020), .ZN(n2385) );
  INV_X4 U2274 ( .A(n1330), .ZN(n2341) );
  INV_X4 U2275 ( .A(n1320), .ZN(n2342) );
  NOR2_X2 U2276 ( .A1(n1551), .A2(n364), .ZN(n1320) );
  INV_X4 U2277 ( .A(n2020), .ZN(n2387) );
  INV_X4 U2278 ( .A(n978), .ZN(n2438) );
  NAND3_X2 U2279 ( .A1(n2433), .A2(n2428), .A3(n719), .ZN(n634) );
  NAND3_X2 U2280 ( .A1(n2433), .A2(n2428), .A3(n719), .ZN(n2337) );
  NAND3_X2 U2281 ( .A1(n2433), .A2(n2428), .A3(n719), .ZN(n2336) );
  INV_X4 U2282 ( .A(n2423), .ZN(n2422) );
  INV_X4 U2283 ( .A(n2360), .ZN(n2363) );
  INV_X4 U2284 ( .A(n2428), .ZN(n2426) );
  INV_X4 U2285 ( .A(n2321), .ZN(n2352) );
  INV_X4 U2286 ( .A(n2321), .ZN(n2351) );
  INV_X4 U2287 ( .A(n2318), .ZN(n2401) );
  INV_X4 U2288 ( .A(n2318), .ZN(n2402) );
  INV_X4 U2289 ( .A(n2419), .ZN(n2416) );
  INV_X4 U2290 ( .A(n2418), .ZN(n2415) );
  INV_X4 U2291 ( .A(n2433), .ZN(n2431) );
  INV_X4 U2292 ( .A(n2433), .ZN(n2430) );
  INV_X4 U2293 ( .A(n2419), .ZN(n2417) );
  INV_X4 U2294 ( .A(n2433), .ZN(n2432) );
  INV_X4 U2295 ( .A(n2413), .ZN(n2414) );
  INV_X4 U2296 ( .A(n2024), .ZN(n2338) );
  NOR2_X2 U2297 ( .A1(n405), .A2(n719), .ZN(n641) );
  INV_X4 U2298 ( .A(n2318), .ZN(n2403) );
  INV_X4 U2299 ( .A(n2319), .ZN(n2410) );
  INV_X4 U2300 ( .A(n2319), .ZN(n2411) );
  INV_X4 U2301 ( .A(n2320), .ZN(n2368) );
  INV_X4 U2302 ( .A(n2320), .ZN(n2367) );
  INV_X4 U2303 ( .A(n2319), .ZN(n2412) );
  INV_X4 U2304 ( .A(n2321), .ZN(n2353) );
  INV_X4 U2305 ( .A(n2320), .ZN(n2369) );
  INV_X4 U2306 ( .A(n2017), .ZN(n2407) );
  INV_X4 U2307 ( .A(n2017), .ZN(n2408) );
  INV_X4 U2308 ( .A(n2017), .ZN(n2409) );
  INV_X4 U2309 ( .A(n2428), .ZN(n2427) );
  INV_X4 U2310 ( .A(n2396), .ZN(n2395) );
  AOI21_X2 U2311 ( .B1(n761), .B2(n2444), .A(n773), .ZN(n762) );
  AOI222_X1 U2312 ( .A1(n2314), .A2(n369), .B1(n1575), .B2(n368), .C1(n371), 
        .C2(n2380), .ZN(n1574) );
  AOI222_X1 U2313 ( .A1(n2380), .A2(n368), .B1(n351), .B2(n1575), .C1(n371), 
        .C2(n2314), .ZN(n1573) );
  NOR2_X2 U2314 ( .A1(n1117), .A2(n1114), .ZN(n1575) );
  OAI21_X2 U2315 ( .B1(n974), .B2(n1552), .A(n1579), .ZN(n1551) );
  NAND3_X2 U2316 ( .A1(n1552), .A2(n2383), .A3(n366), .ZN(n1579) );
  NAND3_X2 U2317 ( .A1(n1403), .A2(n1443), .A3(n508), .ZN(n1442) );
  AOI21_X2 U2318 ( .B1(n1494), .B2(n1405), .A(n1495), .ZN(n1493) );
  NAND3_X2 U2319 ( .A1(n1403), .A2(n1337), .A3(n1494), .ZN(n1492) );
  NOR2_X2 U2320 ( .A1(n1491), .A2(n1444), .ZN(n1494) );
  AOI21_X2 U2321 ( .B1(n1469), .B2(n1604), .A(n273), .ZN(n1315) );
  AOI21_X2 U2322 ( .B1(n481), .B2(n1443), .A(n1445), .ZN(n1362) );
  AOI21_X2 U2323 ( .B1(n891), .B2(n2444), .A(n773), .ZN(n892) );
  AOI21_X2 U2324 ( .B1(n884), .B2(n2444), .A(n773), .ZN(n885) );
  AOI21_X2 U2325 ( .B1(n877), .B2(n2444), .A(n773), .ZN(n878) );
  AOI21_X2 U2326 ( .B1(n869), .B2(n2444), .A(n773), .ZN(n871) );
  AOI21_X2 U2327 ( .B1(n850), .B2(n2444), .A(n773), .ZN(n863) );
  AOI21_X2 U2328 ( .B1(n836), .B2(n2444), .A(n773), .ZN(n837) );
  AOI21_X2 U2329 ( .B1(n829), .B2(n2444), .A(n773), .ZN(n830) );
  AOI21_X2 U2330 ( .B1(n822), .B2(n2443), .A(n773), .ZN(n823) );
  AOI21_X2 U2331 ( .B1(n815), .B2(n2444), .A(n773), .ZN(n816) );
  AOI21_X2 U2332 ( .B1(n1471), .B2(n1424), .A(n1462), .ZN(n1423) );
  OAI21_X2 U2333 ( .B1(n1505), .B2(n1506), .A(n1496), .ZN(n1445) );
  NOR2_X2 U2334 ( .A1(n1503), .A2(n1315), .ZN(n1443) );
  NAND3_X2 U2335 ( .A1(n1425), .A2(n1322), .A3(n1465), .ZN(n1386) );
  OAI21_X2 U2336 ( .B1(n1496), .B2(n1497), .A(n1498), .ZN(n1405) );
  AOI21_X2 U2337 ( .B1(n1470), .B2(n1425), .A(n1471), .ZN(n1385) );
  AOI21_X2 U2338 ( .B1(n262), .B2(n1465), .A(n1470), .ZN(n1420) );
  NOR2_X2 U2339 ( .A1(n2373), .A2(n297), .ZN(n618) );
  OAI21_X2 U2340 ( .B1(n1504), .B2(n1503), .A(n1505), .ZN(n1402) );
  NAND3_X2 U2341 ( .A1(n1118), .A2(n974), .A3(n366), .ZN(n1116) );
  NAND3_X2 U2342 ( .A1(n1468), .A2(n277), .A3(n1469), .ZN(n1467) );
  INV_X4 U2343 ( .A(n2323), .ZN(n2383) );
  NOR2_X2 U2344 ( .A1(n1423), .A2(n956), .ZN(n1526) );
  OAI21_X2 U2345 ( .B1(n1498), .B2(n1444), .A(n1490), .ZN(n1564) );
  INV_X4 U2346 ( .A(n2323), .ZN(n2384) );
  NOR2_X2 U2347 ( .A1(n977), .A2(n2426), .ZN(n967) );
  NOR2_X2 U2348 ( .A1(n1850), .A2(n719), .ZN(n639) );
  OAI21_X2 U2349 ( .B1(n666), .B2(n667), .A(n668), .ZN(n633) );
  OR2_X2 U2350 ( .A1(n915), .A2(n2017), .ZN(n2318) );
  OAI21_X2 U2351 ( .B1(n610), .B2(n41), .A(n581), .ZN(n583) );
  NOR2_X2 U2352 ( .A1(n1497), .A2(n1506), .ZN(n1403) );
  NOR3_X2 U2353 ( .A1(n528), .A2(n953), .A3(n956), .ZN(n951) );
  AOI21_X2 U2354 ( .B1(n413), .B2(n681), .A(n61), .ZN(n713) );
  AOI21_X2 U2355 ( .B1(n801), .B2(n2443), .A(n773), .ZN(n802) );
  AOI21_X2 U2356 ( .B1(n808), .B2(n2444), .A(n773), .ZN(n809) );
  AOI21_X2 U2357 ( .B1(n794), .B2(n2444), .A(n773), .ZN(n795) );
  INV_X4 U2358 ( .A(n1844), .ZN(n438) );
  AOI21_X2 U2359 ( .B1(n1462), .B2(n1463), .A(n1464), .ZN(n954) );
  NOR2_X2 U2360 ( .A1(n69), .A2(n915), .ZN(n610) );
  OAI21_X2 U2361 ( .B1(n1685), .B2(n2363), .A(n2340), .ZN(n1691) );
  OAI21_X2 U2362 ( .B1(n443), .B2(n63), .A(n678), .ZN(n691) );
  AND2_X2 U2363 ( .A1(n103), .A2(n2407), .ZN(n2319) );
  AND2_X2 U2364 ( .A1(n120), .A2(n104), .ZN(n2320) );
  INV_X4 U2365 ( .A(n2023), .ZN(n2433) );
  INV_X4 U2366 ( .A(n631), .ZN(n2428) );
  NOR2_X2 U2367 ( .A1(n961), .A2(n953), .ZN(n959) );
  OR2_X2 U2368 ( .A1(n2414), .A2(n120), .ZN(n2321) );
  INV_X4 U2369 ( .A(n2327), .ZN(n2418) );
  INV_X4 U2370 ( .A(n719), .ZN(n2424) );
  INV_X4 U2371 ( .A(n901), .ZN(n2396) );
  INV_X4 U2372 ( .A(n2325), .ZN(n2398) );
  INV_X4 U2373 ( .A(n2325), .ZN(n2399) );
  INV_X4 U2374 ( .A(n2023), .ZN(n2435) );
  INV_X4 U2375 ( .A(n2329), .ZN(n2404) );
  INV_X4 U2376 ( .A(n2023), .ZN(n2434) );
  INV_X4 U2377 ( .A(n719), .ZN(n2423) );
  INV_X4 U2378 ( .A(n2329), .ZN(n2405) );
  INV_X4 U2379 ( .A(n2361), .ZN(n2360) );
  INV_X4 U2380 ( .A(n1658), .ZN(n2361) );
  NOR2_X2 U2381 ( .A1(n1816), .A2(n899), .ZN(n1658) );
  INV_X4 U2382 ( .A(n2328), .ZN(n2349) );
  INV_X4 U2383 ( .A(n2328), .ZN(n2348) );
  OR2_X2 U2384 ( .A1(n899), .A2(n898), .ZN(n2322) );
  INV_X4 U2385 ( .A(n2327), .ZN(n2419) );
  INV_X4 U2386 ( .A(n2026), .ZN(n2340) );
  INV_X4 U2387 ( .A(n2025), .ZN(n2339) );
  INV_X4 U2388 ( .A(n2325), .ZN(n2400) );
  INV_X4 U2389 ( .A(n2329), .ZN(n2406) );
  INV_X4 U2390 ( .A(n2326), .ZN(n2364) );
  INV_X4 U2391 ( .A(n2326), .ZN(n2365) );
  INV_X4 U2392 ( .A(n2331), .ZN(n2357) );
  INV_X4 U2393 ( .A(n2331), .ZN(n2358) );
  INV_X4 U2394 ( .A(n2330), .ZN(n2354) );
  INV_X4 U2395 ( .A(n2330), .ZN(n2355) );
  INV_X4 U2396 ( .A(n2328), .ZN(n2350) );
  INV_X4 U2397 ( .A(n2326), .ZN(n2366) );
  INV_X4 U2398 ( .A(n2016), .ZN(n2346) );
  INV_X4 U2399 ( .A(n2016), .ZN(n2347) );
  INV_X4 U2400 ( .A(n2018), .ZN(n2345) );
  INV_X4 U2401 ( .A(n2018), .ZN(n2344) );
  INV_X4 U2402 ( .A(n2331), .ZN(n2359) );
  INV_X4 U2403 ( .A(n2330), .ZN(n2356) );
  INV_X4 U2404 ( .A(n901), .ZN(n2397) );
  INV_X4 U2405 ( .A(n719), .ZN(n2425) );
  INV_X4 U2406 ( .A(n631), .ZN(n2429) );
  AOI21_X2 U2407 ( .B1(n1410), .B2(n1411), .A(n1419), .ZN(n1417) );
  AOI222_X1 U2408 ( .A1(n2380), .A2(n351), .B1(n1575), .B2(n1577), .C1(n368), 
        .C2(n2314), .ZN(n1570) );
  AOI21_X2 U2409 ( .B1(n960), .B2(n1543), .A(n1560), .ZN(n1559) );
  NOR3_X2 U2410 ( .A1(n215), .A2(n216), .A3(n217), .ZN(n1685) );
  NOR2_X2 U2411 ( .A1(n1598), .A2(n1601), .ZN(n1469) );
  NOR2_X2 U2412 ( .A1(n1316), .A2(n1314), .ZN(n1468) );
  AOI21_X2 U2413 ( .B1(n1452), .B2(n1451), .A(n1460), .ZN(n1459) );
  OAI21_X2 U2414 ( .B1(n1514), .B2(n1515), .A(n1523), .ZN(n1521) );
  OAI21_X2 U2415 ( .B1(n250), .B2(n1479), .A(n1489), .ZN(n1487) );
  AOI21_X2 U2416 ( .B1(n1549), .B2(n962), .A(n957), .ZN(n1557) );
  AOI21_X2 U2417 ( .B1(n1376), .B2(n955), .A(n1384), .ZN(n1383) );
  AOI21_X2 U2418 ( .B1(n1432), .B2(n1431), .A(n1440), .ZN(n1439) );
  NAND3_X2 U2419 ( .A1(n1323), .A2(n1328), .A3(n1468), .ZN(n1503) );
  AOI21_X2 U2420 ( .B1(n1603), .B2(n1469), .A(n1539), .ZN(n1504) );
  NAND3_X2 U2421 ( .A1(n1393), .A2(n504), .A3(n1400), .ZN(n1531) );
  AOI21_X2 U2422 ( .B1(n187), .B2(n2362), .A(n1796), .ZN(n1801) );
  AOI21_X2 U2423 ( .B1(n220), .B2(n2362), .A(n1781), .ZN(n1786) );
  NAND3_X2 U2424 ( .A1(n1452), .A2(n516), .A3(n1458), .ZN(n1561) );
  AOI21_X2 U2425 ( .B1(n1539), .B2(n1468), .A(n1540), .ZN(n1466) );
  NAND3_X2 U2426 ( .A1(n1328), .A2(n1540), .A3(n1323), .ZN(n1563) );
  NAND3_X2 U2427 ( .A1(n1376), .A2(n1535), .A3(n1382), .ZN(n1566) );
  NAND3_X2 U2428 ( .A1(n976), .A2(n2020), .A3(n1589), .ZN(n978) );
  NOR2_X2 U2429 ( .A1(n1597), .A2(n1502), .ZN(n1604) );
  OAI21_X2 U2430 ( .B1(n1776), .B2(n2361), .A(n2340), .ZN(n1781) );
  OAI21_X2 U2431 ( .B1(n1806), .B2(n2363), .A(n2340), .ZN(n1811) );
  OAI21_X2 U2432 ( .B1(n1791), .B2(n2361), .A(n2340), .ZN(n1796) );
  OAI21_X2 U2433 ( .B1(n1766), .B2(n2361), .A(n2340), .ZN(n1771) );
  OAI21_X2 U2434 ( .B1(n1756), .B2(n2361), .A(n2340), .ZN(n1761) );
  OAI21_X2 U2435 ( .B1(n1746), .B2(n2361), .A(n2340), .ZN(n1751) );
  OAI21_X2 U2436 ( .B1(n1736), .B2(n2363), .A(n2340), .ZN(n1741) );
  OAI21_X2 U2437 ( .B1(n1726), .B2(n2363), .A(n2340), .ZN(n1731) );
  OAI21_X2 U2438 ( .B1(n1716), .B2(n2363), .A(n2340), .ZN(n1721) );
  AOI222_X1 U2439 ( .A1(n370), .A2(n2377), .B1(n373), .B2(n2436), .C1(n535), 
        .C2(n2385), .ZN(n1586) );
  NOR2_X2 U2440 ( .A1(n2381), .A2(n1295), .ZN(n626) );
  NOR2_X2 U2441 ( .A1(n1603), .A2(n1604), .ZN(n1599) );
  NAND3_X2 U2442 ( .A1(n1344), .A2(n485), .A3(n1338), .ZN(n1537) );
  NAND3_X2 U2443 ( .A1(n1411), .A2(n506), .A3(n1418), .ZN(n1565) );
  AOI222_X1 U2444 ( .A1(n372), .A2(n2377), .B1(n374), .B2(n2436), .C1(n370), 
        .C2(n2385), .ZN(n1588) );
  OAI21_X2 U2445 ( .B1(n1392), .B2(n509), .A(n1401), .ZN(n1399) );
  NOR2_X2 U2446 ( .A1(n1501), .A2(n1502), .ZN(n1499) );
  AOI222_X1 U2447 ( .A1(n535), .A2(n2377), .B1(n372), .B2(n2436), .C1(n384), 
        .C2(n2385), .ZN(n1581) );
  NOR2_X2 U2448 ( .A1(n2324), .A2(n974), .ZN(n2323) );
  XNOR2_X2 U2449 ( .A(n376), .B(n2019), .ZN(n2324) );
  AOI222_X1 U2450 ( .A1(n384), .A2(n2377), .B1(n370), .B2(n2436), .C1(n534), 
        .C2(n2385), .ZN(n1576) );
  AOI21_X2 U2451 ( .B1(n1839), .B2(n650), .A(n694), .ZN(n1883) );
  AOI21_X2 U2452 ( .B1(n1839), .B2(n440), .A(n694), .ZN(n1891) );
  AOI21_X2 U2453 ( .B1(n1839), .B2(n670), .A(n694), .ZN(n1897) );
  AOI222_X1 U2454 ( .A1(n456), .A2(n2018), .B1(n457), .B2(n2016), .C1(n455), 
        .C2(n441), .ZN(n686) );
  NOR2_X2 U2455 ( .A1(n718), .A2(n719), .ZN(n681) );
  AOI21_X2 U2456 ( .B1(n638), .B2(n1839), .A(n694), .ZN(n1879) );
  AOI21_X2 U2457 ( .B1(n1337), .B2(n1338), .A(n1345), .ZN(n1343) );
  AOI21_X2 U2458 ( .B1(n1322), .B2(n1323), .A(n1329), .ZN(n1327) );
  OAI21_X2 U2459 ( .B1(n612), .B2(n169), .A(n901), .ZN(n1592) );
  OR2_X2 U2460 ( .A1(n611), .A2(n2017), .ZN(n2325) );
  OAI21_X2 U2461 ( .B1(n42), .B2(n2423), .A(n455), .ZN(n720) );
  NOR2_X2 U2462 ( .A1(n672), .A2(n666), .ZN(n637) );
  OAI21_X2 U2463 ( .B1(n1315), .B2(n1316), .A(n1317), .ZN(n1313) );
  AOI21_X2 U2464 ( .B1(n402), .B2(n712), .A(n400), .ZN(n1911) );
  NOR2_X2 U2465 ( .A1(n1479), .A2(n1488), .ZN(n1542) );
  NAND3_X2 U2466 ( .A1(n454), .A2(n397), .A3(n101), .ZN(n1649) );
  NAND3_X2 U2467 ( .A1(n1458), .A2(n1452), .A3(n1542), .ZN(n956) );
  OAI21_X2 U2468 ( .B1(n1638), .B2(n1644), .A(n2393), .ZN(n1611) );
  OAI21_X2 U2469 ( .B1(n1638), .B2(n1641), .A(n2392), .ZN(n1608) );
  OAI21_X2 U2470 ( .B1(n1638), .B2(n1642), .A(n2392), .ZN(n1609) );
  OAI21_X2 U2471 ( .B1(n1638), .B2(n1643), .A(n2392), .ZN(n1610) );
  OAI21_X2 U2472 ( .B1(n1638), .B2(n1645), .A(n2392), .ZN(n1612) );
  OAI21_X2 U2473 ( .B1(n1638), .B2(n1646), .A(n2392), .ZN(n1613) );
  OAI21_X2 U2474 ( .B1(n1638), .B2(n1639), .A(n2392), .ZN(n1605) );
  OAI21_X2 U2475 ( .B1(n1638), .B2(n1640), .A(n2392), .ZN(n1607) );
  OAI21_X2 U2476 ( .B1(n1639), .B2(n1648), .A(n2393), .ZN(n1622) );
  OAI21_X2 U2477 ( .B1(n1640), .B2(n1648), .A(n2393), .ZN(n1623) );
  OAI21_X2 U2478 ( .B1(n1641), .B2(n1648), .A(n2393), .ZN(n1624) );
  OAI21_X2 U2479 ( .B1(n1642), .B2(n1648), .A(n2393), .ZN(n1625) );
  OAI21_X2 U2480 ( .B1(n1643), .B2(n1648), .A(n2393), .ZN(n1626) );
  OAI21_X2 U2481 ( .B1(n1644), .B2(n1648), .A(n2393), .ZN(n1627) );
  OAI21_X2 U2482 ( .B1(n1645), .B2(n1648), .A(n2393), .ZN(n1628) );
  OAI21_X2 U2483 ( .B1(n1646), .B2(n1648), .A(n2394), .ZN(n1629) );
  AOI21_X2 U2484 ( .B1(n398), .B2(n2443), .A(n773), .ZN(n777) );
  OAI21_X2 U2485 ( .B1(n1643), .B2(n1647), .A(n2393), .ZN(n1618) );
  OAI21_X2 U2486 ( .B1(n1644), .B2(n1647), .A(n2393), .ZN(n1619) );
  OAI21_X2 U2487 ( .B1(n1645), .B2(n1647), .A(n2393), .ZN(n1620) );
  OAI21_X2 U2488 ( .B1(n1646), .B2(n1647), .A(n2393), .ZN(n1621) );
  OAI21_X2 U2489 ( .B1(n1639), .B2(n1647), .A(n2392), .ZN(n1614) );
  OAI21_X2 U2490 ( .B1(n1640), .B2(n1647), .A(n2392), .ZN(n1615) );
  OAI21_X2 U2491 ( .B1(n1641), .B2(n1647), .A(n2392), .ZN(n1616) );
  OAI21_X2 U2492 ( .B1(n1642), .B2(n1647), .A(n2392), .ZN(n1617) );
  OAI21_X2 U2493 ( .B1(n1639), .B2(n1649), .A(n2394), .ZN(n1630) );
  OAI21_X2 U2494 ( .B1(n1640), .B2(n1649), .A(n2394), .ZN(n1631) );
  OAI21_X2 U2495 ( .B1(n1641), .B2(n1649), .A(n2394), .ZN(n1632) );
  OAI21_X2 U2496 ( .B1(n1643), .B2(n1649), .A(n2394), .ZN(n1634) );
  OAI21_X2 U2497 ( .B1(n1642), .B2(n1649), .A(n2394), .ZN(n1633) );
  OAI21_X2 U2498 ( .B1(n1644), .B2(n1649), .A(n2394), .ZN(n1635) );
  OAI21_X2 U2499 ( .B1(n1645), .B2(n1649), .A(n2392), .ZN(n1636) );
  AOI21_X2 U2500 ( .B1(n786), .B2(n2443), .A(n773), .ZN(n784) );
  INV_X4 U2501 ( .A(n1843), .ZN(n439) );
  NAND3_X2 U2502 ( .A1(n1650), .A2(n1820), .A3(n1819), .ZN(n898) );
  NAND3_X2 U2503 ( .A1(n2419), .A2(n109), .A3(n1653), .ZN(n1652) );
  OAI21_X2 U2504 ( .B1(n107), .B2(n120), .A(n898), .ZN(n1653) );
  NAND3_X2 U2505 ( .A1(n718), .A2(n455), .A3(n2423), .ZN(n678) );
  OAI21_X2 U2506 ( .B1(n1675), .B2(n2361), .A(n2340), .ZN(n1680) );
  OAI21_X2 U2507 ( .B1(n2361), .B2(n399), .A(n2340), .ZN(n1668) );
  NOR2_X2 U2508 ( .A1(n1515), .A2(n1522), .ZN(n960) );
  AOI21_X2 U2509 ( .B1(n520), .B2(n1542), .A(n1543), .ZN(n961) );
  NAND3_X2 U2510 ( .A1(n1819), .A2(n1820), .A3(n120), .ZN(n1816) );
  NAND3_X2 U2511 ( .A1(n1432), .A2(n512), .A3(n1438), .ZN(n1528) );
  NOR2_X2 U2512 ( .A1(n1836), .A2(n718), .ZN(n1872) );
  OAI21_X2 U2513 ( .B1(n1696), .B2(n2363), .A(n2340), .ZN(n1701) );
  OAI21_X2 U2514 ( .B1(n1706), .B2(n2363), .A(n2340), .ZN(n1711) );
  AOI21_X2 U2515 ( .B1(n1349), .B2(n1350), .A(n1356), .ZN(n1354) );
  NOR2_X2 U2516 ( .A1(n298), .A2(n2020), .ZN(n624) );
  NAND3_X2 U2517 ( .A1(n393), .A2(n394), .A3(n396), .ZN(n1646) );
  INV_X4 U2518 ( .A(n756), .ZN(n40) );
  NOR3_X2 U2519 ( .A1(n217), .A2(n216), .A3(n2363), .ZN(n1681) );
  NAND3_X2 U2520 ( .A1(n585), .A2(n584), .A3(n595), .ZN(n600) );
  OAI21_X2 U2521 ( .B1(n1599), .B2(n1598), .A(n1602), .ZN(n1600) );
  OAI21_X2 U2522 ( .B1(n1362), .B2(n494), .A(n1370), .ZN(n1368) );
  NAND3_X2 U2523 ( .A1(n2418), .A2(n109), .A3(n106), .ZN(n899) );
  NAND3_X2 U2524 ( .A1(n968), .A2(n479), .A3(n104), .ZN(n613) );
  AND2_X2 U2525 ( .A1(n104), .A2(n1650), .ZN(n2326) );
  AND2_X2 U2526 ( .A1(n612), .A2(n2433), .ZN(n2327) );
  AOI21_X2 U2527 ( .B1(n681), .B2(n712), .A(n61), .ZN(n711) );
  OR2_X2 U2528 ( .A1(n1650), .A2(n2414), .ZN(n2328) );
  OR2_X2 U2529 ( .A1(n916), .A2(n2017), .ZN(n2329) );
  OR2_X2 U2530 ( .A1(n898), .A2(n2333), .ZN(n2330) );
  OR2_X2 U2531 ( .A1(n1816), .A2(n2333), .ZN(n2331) );
  INV_X4 U2532 ( .A(n2333), .ZN(n2420) );
  INV_X4 U2533 ( .A(n2332), .ZN(n2393) );
  INV_X4 U2534 ( .A(n2332), .ZN(n2392) );
  INV_X4 U2535 ( .A(n2333), .ZN(n2421) );
  INV_X4 U2536 ( .A(n2332), .ZN(n2394) );
  INV_X4 U2537 ( .A(n757), .ZN(n2413) );
  NOR2_X2 U2538 ( .A1(n916), .A2(n69), .ZN(n631) );
  AOI21_X2 U2539 ( .B1(n216), .B2(n2362), .A(n1680), .ZN(n1686) );
  OAI21_X2 U2540 ( .B1(q[29]), .B2(n2322), .A(n762), .ZN(n759) );
  NOR3_X2 U2541 ( .A1(n761), .A2(q[29]), .A3(n2441), .ZN(n897) );
  NAND3_X2 U2542 ( .A1(q[1]), .A2(q[0]), .A3(q[2]), .ZN(n786) );
  AOI222_X1 U2543 ( .A1(n2375), .A2(sdata[25]), .B1(n2436), .B2(sdata[23]), 
        .C1(n2387), .C2(sdata[26]), .ZN(n1577) );
  AOI222_X1 U2544 ( .A1(n2376), .A2(sdata[6]), .B1(n2438), .B2(sdata[4]), .C1(
        n2385), .C2(sdata[7]), .ZN(n1374) );
  AOI222_X1 U2545 ( .A1(n2376), .A2(sdata[7]), .B1(n2438), .B2(sdata[5]), .C1(
        n2386), .C2(sdata[8]), .ZN(n1380) );
  AOI222_X1 U2546 ( .A1(n2376), .A2(sdata[8]), .B1(n2438), .B2(sdata[6]), .C1(
        n2385), .C2(sdata[9]), .ZN(n1390) );
  AOI222_X1 U2547 ( .A1(n2375), .A2(sdata[19]), .B1(n2437), .B2(sdata[17]), 
        .C1(n2386), .C2(sdata[20]), .ZN(n1519) );
  AOI222_X1 U2548 ( .A1(n2375), .A2(sdata[17]), .B1(n2437), .B2(sdata[15]), 
        .C1(n2386), .C2(sdata[18]), .ZN(n1484) );
  AOI222_X1 U2549 ( .A1(n2375), .A2(sdata[21]), .B1(n2436), .B2(sdata[19]), 
        .C1(n2386), .C2(sdata[22]), .ZN(n1554) );
  AOI222_X1 U2550 ( .A1(n2376), .A2(sdata[5]), .B1(n2437), .B2(sdata[3]), .C1(
        n2385), .C2(sdata[6]), .ZN(n1366) );
  AOI222_X1 U2551 ( .A1(n2376), .A2(sdata[9]), .B1(n2437), .B2(sdata[7]), .C1(
        n2385), .C2(sdata[10]), .ZN(n1397) );
  AOI222_X1 U2552 ( .A1(n2376), .A2(sdata[10]), .B1(n2437), .B2(sdata[8]), 
        .C1(n2385), .C2(sdata[11]), .ZN(n1408) );
  AOI222_X1 U2553 ( .A1(n2376), .A2(sdata[11]), .B1(n2437), .B2(sdata[9]), 
        .C1(n2386), .C2(sdata[12]), .ZN(n1414) );
  AOI222_X1 U2554 ( .A1(n2376), .A2(sdata[12]), .B1(n2437), .B2(sdata[10]), 
        .C1(n2386), .C2(sdata[13]), .ZN(n1428) );
  AOI222_X1 U2555 ( .A1(n2375), .A2(sdata[20]), .B1(n2436), .B2(sdata[18]), 
        .C1(n2386), .C2(sdata[21]), .ZN(n1547) );
  AOI222_X1 U2556 ( .A1(n2376), .A2(sdata[4]), .B1(n2436), .B2(sdata[2]), .C1(
        n2385), .C2(sdata[5]), .ZN(n1360) );
  AOI222_X1 U2557 ( .A1(n2375), .A2(sdata[14]), .B1(n2437), .B2(sdata[12]), 
        .C1(n2386), .C2(sdata[15]), .ZN(n1448) );
  AOI222_X1 U2558 ( .A1(n2375), .A2(sdata[16]), .B1(n2437), .B2(sdata[14]), 
        .C1(n2386), .C2(sdata[17]), .ZN(n1475) );
  AOI222_X1 U2559 ( .A1(n2375), .A2(sdata[18]), .B1(n2437), .B2(sdata[16]), 
        .C1(n2386), .C2(sdata[19]), .ZN(n1511) );
  AOI222_X1 U2560 ( .A1(n2375), .A2(sdata[22]), .B1(n2437), .B2(sdata[20]), 
        .C1(n2387), .C2(sdata[23]), .ZN(n1571) );
  AOI222_X1 U2561 ( .A1(n2376), .A2(sdata[13]), .B1(n2437), .B2(sdata[11]), 
        .C1(n2386), .C2(sdata[14]), .ZN(n1435) );
  AOI222_X1 U2562 ( .A1(n2375), .A2(sdata[15]), .B1(n2437), .B2(sdata[13]), 
        .C1(n2386), .C2(sdata[16]), .ZN(n1455) );
  AOI222_X1 U2563 ( .A1(n2375), .A2(sdata[24]), .B1(n2436), .B2(sdata[22]), 
        .C1(n2386), .C2(sdata[25]), .ZN(n1578) );
  AOI222_X1 U2564 ( .A1(n2375), .A2(sdata[23]), .B1(n2436), .B2(sdata[21]), 
        .C1(n2387), .C2(sdata[24]), .ZN(n1572) );
  AOI222_X1 U2565 ( .A1(n2376), .A2(sdata[3]), .B1(sdata[1]), .B2(n2436), .C1(
        n2385), .C2(sdata[4]), .ZN(n1335) );
  AOI222_X1 U2566 ( .A1(n2376), .A2(sdata[2]), .B1(sdata[0]), .B2(n2436), .C1(
        n2385), .C2(sdata[3]), .ZN(n1308) );
  NAND3_X2 U2567 ( .A1(n942), .A2(n943), .A3(n950), .ZN(n933) );
  OAI21_X2 U2568 ( .B1(q[25]), .B2(n2442), .A(n885), .ZN(n887) );
  OAI21_X2 U2569 ( .B1(q[23]), .B2(n2441), .A(n878), .ZN(n880) );
  NOR3_X2 U2570 ( .A1(n2441), .A2(q[27]), .A3(n891), .ZN(n890) );
  OAI21_X2 U2571 ( .B1(q[21]), .B2(n2442), .A(n871), .ZN(n873) );
  OAI21_X2 U2572 ( .B1(q[19]), .B2(n2442), .A(n863), .ZN(n865) );
  OAI21_X2 U2573 ( .B1(q[17]), .B2(n2442), .A(n837), .ZN(n842) );
  NOR3_X2 U2574 ( .A1(n2441), .A2(q[25]), .A3(n884), .ZN(n883) );
  NOR3_X2 U2575 ( .A1(n2441), .A2(q[21]), .A3(n869), .ZN(n868) );
  OAI21_X2 U2576 ( .B1(q[27]), .B2(n2322), .A(n892), .ZN(n894) );
  OAI21_X2 U2577 ( .B1(q[15]), .B2(n2322), .A(n830), .ZN(n832) );
  OAI21_X2 U2578 ( .B1(q[13]), .B2(n2322), .A(n823), .ZN(n825) );
  OAI21_X2 U2579 ( .B1(q[11]), .B2(n2322), .A(n816), .ZN(n818) );
  AOI222_X1 U2580 ( .A1(n2404), .A2(i_dividend[31]), .B1(n2403), .B2(n2019), 
        .C1(n2400), .C2(n769), .ZN(n765) );
  AOI222_X1 U2581 ( .A1(n2405), .A2(i_dividend[28]), .B1(n2401), .B2(n330), 
        .C1(n930), .C2(n2398), .ZN(n1520) );
  AOI222_X1 U2582 ( .A1(n2404), .A2(i_dividend[30]), .B1(n2401), .B2(n346), 
        .C1(n932), .C2(n2398), .ZN(n1556) );
  AOI222_X1 U2583 ( .A1(i_dividend[2]), .A2(n2406), .B1(n2403), .B2(n615), 
        .C1(n1299), .C2(n2400), .ZN(n1298) );
  AOI222_X1 U2584 ( .A1(i_dividend[7]), .A2(n2405), .B1(n2402), .B2(n291), 
        .C1(n269), .C2(n2399), .ZN(n1321) );
  AOI222_X1 U2585 ( .A1(i_dividend[6]), .A2(n2406), .B1(n2403), .B2(n292), 
        .C1(n917), .C2(n2400), .ZN(n1312) );
  AOI222_X1 U2586 ( .A1(i_dividend[3]), .A2(n2406), .B1(n2403), .B2(n618), 
        .C1(n276), .C2(n2400), .ZN(n1303) );
  AOI222_X1 U2587 ( .A1(i_dividend[4]), .A2(n2406), .B1(n2403), .B2(n620), 
        .C1(n275), .C2(n2400), .ZN(n1305) );
  AOI222_X1 U2588 ( .A1(i_dividend[5]), .A2(n2406), .B1(n2403), .B2(n622), 
        .C1(n1310), .C2(n2400), .ZN(n1309) );
  AOI222_X1 U2589 ( .A1(n2405), .A2(i_dividend[29]), .B1(n2401), .B2(n347), 
        .C1(n931), .C2(n2398), .ZN(n1548) );
  AOI222_X1 U2590 ( .A1(n2404), .A2(i_dividend[18]), .B1(n2402), .B2(n736), 
        .C1(n923), .C2(n2399), .ZN(n1398) );
  AOI222_X1 U2591 ( .A1(n2405), .A2(i_dividend[21]), .B1(n2401), .B2(n740), 
        .C1(n924), .C2(n2398), .ZN(n1430) );
  AOI222_X1 U2592 ( .A1(n2405), .A2(i_dividend[23]), .B1(n2401), .B2(n743), 
        .C1(n926), .C2(n2398), .ZN(n1450) );
  AOI222_X1 U2593 ( .A1(n2405), .A2(i_dividend[24]), .B1(n2401), .B2(n745), 
        .C1(n927), .C2(n2398), .ZN(n1457) );
  AOI222_X1 U2594 ( .A1(n2405), .A2(i_dividend[26]), .B1(n2401), .B2(n748), 
        .C1(n928), .C2(n2398), .ZN(n1486) );
  AOI222_X1 U2595 ( .A1(n2405), .A2(i_dividend[27]), .B1(n2401), .B2(n750), 
        .C1(n929), .C2(n2398), .ZN(n1513) );
  AOI222_X1 U2596 ( .A1(i_dividend[1]), .A2(n2406), .B1(n2403), .B2(n626), 
        .C1(n1123), .C2(n2400), .ZN(n1122) );
  NOR3_X2 U2597 ( .A1(n2441), .A2(q[15]), .A3(n829), .ZN(n828) );
  AOI222_X1 U2598 ( .A1(n2405), .A2(i_dividend[25]), .B1(n2401), .B2(n746), 
        .C1(n251), .C2(n2398), .ZN(n1477) );
  AOI222_X1 U2599 ( .A1(n2404), .A2(i_dividend[19]), .B1(n2401), .B2(n737), 
        .C1(n261), .C2(n2398), .ZN(n1409) );
  AOI222_X1 U2600 ( .A1(n2404), .A2(i_dividend[20]), .B1(n2401), .B2(n739), 
        .C1(n260), .C2(n2398), .ZN(n1416) );
  AOI222_X1 U2601 ( .A1(n2405), .A2(i_dividend[22]), .B1(n2401), .B2(n742), 
        .C1(n925), .C2(n2398), .ZN(n1437) );
  AOI21_X2 U2602 ( .B1(n184), .B2(n2362), .A(n1811), .ZN(n1815) );
  NOR3_X2 U2603 ( .A1(n3284), .A2(n3285), .A3(n218), .ZN(n1675) );
  OAI21_X2 U2604 ( .B1(n2387), .B2(n976), .A(n978), .ZN(n972) );
  NAND3_X2 U2605 ( .A1(n1120), .A2(n1118), .A3(n367), .ZN(n1119) );
  AOI222_X1 U2606 ( .A1(reg_a[29]), .A2(n2415), .B1(n2351), .B2(n122), .C1(
        n2348), .C2(n3182), .ZN(n1810) );
  AOI222_X1 U2607 ( .A1(reg_a[26]), .A2(n2415), .B1(n2351), .B2(n125), .C1(
        n2348), .C2(n3176), .ZN(n1795) );
  AOI222_X1 U2608 ( .A1(reg_a[23]), .A2(n2415), .B1(n2351), .B2(n128), .C1(
        n2348), .C2(n3170), .ZN(n1780) );
  AOI222_X1 U2609 ( .A1(reg_a[21]), .A2(n2415), .B1(n2351), .B2(n130), .C1(
        n2348), .C2(n3166), .ZN(n1770) );
  AOI222_X1 U2610 ( .A1(reg_a[19]), .A2(n2416), .B1(n2352), .B2(n132), .C1(
        n2349), .C2(n3162), .ZN(n1760) );
  AOI222_X1 U2611 ( .A1(reg_a[17]), .A2(n2416), .B1(n2352), .B2(n134), .C1(
        n2349), .C2(n3158), .ZN(n1750) );
  AOI222_X1 U2612 ( .A1(reg_a[15]), .A2(n2416), .B1(n2352), .B2(n136), .C1(
        n2349), .C2(n3154), .ZN(n1740) );
  AOI222_X1 U2613 ( .A1(reg_a[13]), .A2(n2416), .B1(n2352), .B2(n138), .C1(
        n2349), .C2(n3150), .ZN(n1730) );
  NOR3_X2 U2614 ( .A1(n2441), .A2(q[23]), .A3(n877), .ZN(n876) );
  NOR3_X2 U2615 ( .A1(n2441), .A2(q[19]), .A3(n850), .ZN(n848) );
  NOR3_X2 U2616 ( .A1(n2441), .A2(q[17]), .A3(n836), .ZN(n835) );
  NOR3_X2 U2617 ( .A1(n2322), .A2(q[13]), .A3(n822), .ZN(n821) );
  NOR3_X2 U2618 ( .A1(n2441), .A2(q[11]), .A3(n815), .ZN(n814) );
  OAI21_X2 U2619 ( .B1(nq[21]), .B2(n2361), .A(n10), .ZN(n1775) );
  OAI21_X2 U2620 ( .B1(nq[19]), .B2(n2361), .A(n11), .ZN(n1765) );
  OAI21_X2 U2621 ( .B1(nq[17]), .B2(n2361), .A(n12), .ZN(n1755) );
  OAI21_X2 U2622 ( .B1(nq[15]), .B2(n2363), .A(n13), .ZN(n1745) );
  OAI21_X2 U2623 ( .B1(nq[13]), .B2(n2363), .A(n14), .ZN(n1735) );
  OAI21_X2 U2624 ( .B1(nq[27]), .B2(n2361), .A(n1801), .ZN(n1805) );
  OAI21_X2 U2625 ( .B1(nq[24]), .B2(n2361), .A(n1786), .ZN(n1790) );
  AOI222_X1 U2626 ( .A1(n2404), .A2(i_dividend[15]), .B1(n2402), .B2(n304), 
        .C1(n921), .C2(n2399), .ZN(n1375) );
  AOI222_X1 U2627 ( .A1(n2404), .A2(i_dividend[17]), .B1(n2402), .B2(n301), 
        .C1(n255), .C2(n2399), .ZN(n1391) );
  AOI222_X1 U2628 ( .A1(n2404), .A2(i_dividend[16]), .B1(n2402), .B2(n302), 
        .C1(n922), .C2(n2399), .ZN(n1381) );
  AOI222_X1 U2629 ( .A1(i_dividend[10]), .A2(n2405), .B1(n2402), .B2(n288), 
        .C1(n252), .C2(n2399), .ZN(n1342) );
  AOI222_X1 U2630 ( .A1(n2404), .A2(i_dividend[12]), .B1(n2402), .B2(n285), 
        .C1(n258), .C2(n2399), .ZN(n1353) );
  AOI222_X1 U2631 ( .A1(n2404), .A2(i_dividend[13]), .B1(n2402), .B2(n307), 
        .C1(n919), .C2(n2399), .ZN(n1361) );
  AOI222_X1 U2632 ( .A1(n2404), .A2(i_dividend[14]), .B1(n2402), .B2(n305), 
        .C1(n920), .C2(n2399), .ZN(n1367) );
  AOI222_X1 U2633 ( .A1(n2404), .A2(i_dividend[11]), .B1(n2402), .B2(n286), 
        .C1(n918), .C2(n2399), .ZN(n1348) );
  NAND3_X2 U2634 ( .A1(n1802), .A2(n1803), .A3(n1804), .ZN(n1014) );
  AOI222_X1 U2635 ( .A1(reg_a[28]), .A2(n2415), .B1(n2351), .B2(n123), .C1(
        n2348), .C2(n3180), .ZN(n1804) );
  NAND3_X2 U2636 ( .A1(n1797), .A2(n1798), .A3(n1799), .ZN(n1015) );
  AOI222_X1 U2637 ( .A1(reg_a[27]), .A2(n2416), .B1(n2351), .B2(n124), .C1(
        n2348), .C2(n3178), .ZN(n1799) );
  NAND3_X2 U2638 ( .A1(n1812), .A2(n7), .A3(n1813), .ZN(n1012) );
  AOI222_X1 U2639 ( .A1(reg_a[30]), .A2(n2415), .B1(n2351), .B2(n121), .C1(
        n2348), .C2(n3184), .ZN(n1813) );
  NAND3_X2 U2640 ( .A1(n1787), .A2(n1788), .A3(n1789), .ZN(n1017) );
  AOI222_X1 U2641 ( .A1(reg_a[25]), .A2(n2415), .B1(n2351), .B2(n126), .C1(
        n2348), .C2(n3174), .ZN(n1789) );
  NAND3_X2 U2642 ( .A1(n1782), .A2(n1783), .A3(n1784), .ZN(n1018) );
  AOI222_X1 U2643 ( .A1(reg_a[24]), .A2(n2415), .B1(n2351), .B2(n127), .C1(
        n2348), .C2(n3172), .ZN(n1784) );
  NAND3_X2 U2644 ( .A1(n1772), .A2(n1773), .A3(n1774), .ZN(n1020) );
  AOI222_X1 U2645 ( .A1(reg_a[22]), .A2(n2415), .B1(n2351), .B2(n129), .C1(
        n2348), .C2(n3168), .ZN(n1774) );
  NAND3_X2 U2646 ( .A1(n1762), .A2(n1763), .A3(n1764), .ZN(n1022) );
  AOI222_X1 U2647 ( .A1(reg_a[20]), .A2(n2416), .B1(n2351), .B2(n131), .C1(
        n2348), .C2(n3164), .ZN(n1764) );
  NAND3_X2 U2648 ( .A1(n1752), .A2(n1753), .A3(n1754), .ZN(n1024) );
  AOI222_X1 U2649 ( .A1(reg_a[18]), .A2(n2416), .B1(n2352), .B2(n133), .C1(
        n2349), .C2(n3160), .ZN(n1754) );
  NAND3_X2 U2650 ( .A1(n1742), .A2(n1743), .A3(n1744), .ZN(n1026) );
  AOI222_X1 U2651 ( .A1(reg_a[16]), .A2(n2416), .B1(n2352), .B2(n135), .C1(
        n2349), .C2(n3156), .ZN(n1744) );
  NAND3_X2 U2652 ( .A1(n1732), .A2(n1733), .A3(n1734), .ZN(n1028) );
  AOI222_X1 U2653 ( .A1(reg_a[14]), .A2(n2416), .B1(n2352), .B2(n137), .C1(
        n2349), .C2(n3152), .ZN(n1734) );
  NAND3_X2 U2654 ( .A1(n1722), .A2(n1723), .A3(n1724), .ZN(n1030) );
  AOI222_X1 U2655 ( .A1(reg_a[12]), .A2(n2416), .B1(n2352), .B2(n139), .C1(
        n2349), .C2(n3148), .ZN(n1724) );
  AOI222_X1 U2656 ( .A1(i_dividend[9]), .A2(n2405), .B1(n2402), .B2(n289), 
        .C1(n253), .C2(n2399), .ZN(n1336) );
  AOI222_X1 U2657 ( .A1(i_dividend[8]), .A2(n2406), .B1(n2402), .B2(n290), 
        .C1(n268), .C2(n2399), .ZN(n1326) );
  NAND3_X2 U2658 ( .A1(n2360), .A2(nq[21]), .A3(n1766), .ZN(n1768) );
  NAND3_X2 U2659 ( .A1(n1658), .A2(nq[19]), .A3(n1756), .ZN(n1758) );
  NAND3_X2 U2660 ( .A1(n1658), .A2(nq[17]), .A3(n1746), .ZN(n1748) );
  NAND3_X2 U2661 ( .A1(n1658), .A2(nq[15]), .A3(n1736), .ZN(n1738) );
  NAND3_X2 U2662 ( .A1(n1658), .A2(nq[13]), .A3(n1726), .ZN(n1728) );
  NAND3_X2 U2663 ( .A1(n2360), .A2(nq[29]), .A3(n1806), .ZN(n1808) );
  NAND3_X2 U2664 ( .A1(n1658), .A2(nq[23]), .A3(n1776), .ZN(n1778) );
  NAND3_X2 U2665 ( .A1(n1658), .A2(nq[26]), .A3(n1791), .ZN(n1793) );
  OAI21_X2 U2666 ( .B1(nq[11]), .B2(n2363), .A(n15), .ZN(n1725) );
  NOR2_X2 U2667 ( .A1(n414), .A2(n946), .ZN(n1839) );
  NOR2_X2 U2668 ( .A1(n1954), .A2(state_reg_1_0), .ZN(n968) );
  AOI222_X1 U2669 ( .A1(reg_b[3]), .A2(n2417), .B1(n2420), .B2(n477), .C1(
        n2413), .C2(n3126), .ZN(n782) );
  AOI222_X1 U2670 ( .A1(n951), .A2(n503), .B1(reg_a[30]), .B2(reg_b[30]), .C1(
        n530), .C2(n952), .ZN(n950) );
  NAND2_X2 U2671 ( .A1(n947), .A2(n946), .ZN(n672) );
  AOI211_X2 U2672 ( .C1(n403), .C2(n1847), .A(n1848), .B(n1849), .ZN(n1845) );
  AOI211_X2 U2673 ( .C1(n1872), .C2(n1873), .A(n1874), .B(n1875), .ZN(n1870)
         );
  AOI211_X2 U2674 ( .C1(n403), .C2(n1861), .A(n1862), .B(n1863), .ZN(n1859) );
  NOR3_X2 U2675 ( .A1(n1937), .A2(n1938), .A3(n1939), .ZN(n1935) );
  NOR3_X2 U2676 ( .A1(n1916), .A2(n1917), .A3(n1918), .ZN(n1914) );
  NOR3_X2 U2677 ( .A1(n1927), .A2(n1928), .A3(n1929), .ZN(n1925) );
  OAI21_X2 U2678 ( .B1(q[9]), .B2(n2322), .A(n809), .ZN(n811) );
  OAI21_X2 U2679 ( .B1(q[5]), .B2(n2322), .A(n795), .ZN(n797) );
  AOI222_X1 U2680 ( .A1(i_dividend[0]), .A2(n2406), .B1(n2403), .B2(n624), 
        .C1(n2400), .C2(n283), .ZN(n1121) );
  NAND2_X2 U2681 ( .A1(n946), .A2(n414), .ZN(n1836) );
  AOI222_X1 U2682 ( .A1(n284), .A2(n2413), .B1(n455), .B2(n2420), .C1(n2415), 
        .C2(reg_b[31]), .ZN(n721) );
  NAND3_X2 U2683 ( .A1(n936), .A2(n454), .A3(n101), .ZN(n1648) );
  AOI222_X1 U2684 ( .A1(reg_a[9]), .A2(n2415), .B1(n2352), .B2(n142), .C1(
        n2349), .C2(n3142), .ZN(n1710) );
  AOI222_X1 U2685 ( .A1(reg_a[5]), .A2(n2417), .B1(n2353), .B2(n113), .C1(
        n2350), .C2(n3134), .ZN(n1690) );
  AOI222_X1 U2686 ( .A1(reg_a[7]), .A2(n2417), .B1(n2353), .B2(n111), .C1(
        n2350), .C2(n3138), .ZN(n1700) );
  OAI21_X2 U2687 ( .B1(n434), .B2(n2025), .A(n678), .ZN(n695) );
  OAI21_X2 U2688 ( .B1(n434), .B2(n63), .A(n678), .ZN(n677) );
  OAI21_X2 U2689 ( .B1(n686), .B2(n63), .A(n678), .ZN(n685) );
  AOI222_X1 U2690 ( .A1(reg_b[2]), .A2(n2417), .B1(n2420), .B2(n473), .C1(
        n2413), .C2(n3123), .ZN(n778) );
  OAI21_X2 U2691 ( .B1(q[1]), .B2(n2322), .A(n777), .ZN(n780) );
  AOI222_X1 U2692 ( .A1(reg_b[4]), .A2(n2416), .B1(n2420), .B2(n472), .C1(
        n2413), .C2(n3129), .ZN(n787) );
  OAI21_X2 U2693 ( .B1(q[3]), .B2(n2322), .A(n784), .ZN(n789) );
  AOI222_X1 U2694 ( .A1(reg_b[5]), .A2(n2417), .B1(n2420), .B2(n471), .C1(
        n2413), .C2(n3132), .ZN(n791) );
  NAND3_X2 U2695 ( .A1(n935), .A2(n936), .A3(n101), .ZN(n1638) );
  NAND3_X2 U2696 ( .A1(n935), .A2(n397), .A3(n101), .ZN(n1647) );
  NAND3_X2 U2697 ( .A1(n938), .A2(n939), .A3(n937), .ZN(n1639) );
  NAND3_X2 U2698 ( .A1(n938), .A2(n394), .A3(n937), .ZN(n1640) );
  NAND3_X2 U2699 ( .A1(n939), .A2(n393), .A3(n937), .ZN(n1641) );
  NAND3_X2 U2700 ( .A1(n939), .A2(n396), .A3(n938), .ZN(n1643) );
  AOI21_X2 U2701 ( .B1(n2362), .B2(n3284), .A(n1668), .ZN(n1674) );
  NOR3_X2 U2702 ( .A1(state[1]), .A2(state[2]), .A3(state[0]), .ZN(n1590) );
  NOR3_X2 U2703 ( .A1(state[4]), .A2(n2022), .A3(state[3]), .ZN(n1651) );
  NOR2_X2 U2704 ( .A1(n936), .A2(n236), .ZN(n606) );
  AOI222_X1 U2705 ( .A1(n2430), .A2(sdata[28]), .B1(n2338), .B2(n650), .C1(n42), .C2(n458), .ZN(n715) );
  AOI222_X1 U2706 ( .A1(n2430), .A2(sdata[27]), .B1(n2338), .B2(n638), .C1(n42), .C2(n459), .ZN(n714) );
  AOI222_X1 U2707 ( .A1(n2430), .A2(sdata[30]), .B1(n2338), .B2(n670), .C1(n42), .C2(n456), .ZN(n717) );
  NOR2_X2 U2708 ( .A1(n946), .A2(n947), .ZN(n1838) );
  AOI222_X1 U2709 ( .A1(n40), .A2(n445), .B1(n2444), .B2(n398), .C1(n773), 
        .C2(q[0]), .ZN(n771) );
  AOI222_X1 U2710 ( .A1(n2430), .A2(sdata[29]), .B1(n2338), .B2(n440), .C1(n42), .C2(n457), .ZN(n716) );
  NOR2_X2 U2711 ( .A1(n946), .A2(n870), .ZN(n712) );
  NAND3_X2 U2712 ( .A1(n393), .A2(n394), .A3(n937), .ZN(n1642) );
  NAND3_X2 U2713 ( .A1(n104), .A2(n968), .A3(n934), .ZN(n754) );
  NAND3_X2 U2714 ( .A1(n396), .A2(n394), .A3(n938), .ZN(n1644) );
  NAND3_X2 U2715 ( .A1(n396), .A2(n393), .A3(n939), .ZN(n1645) );
  AOI21_X2 U2716 ( .B1(n1680), .B2(n216), .A(n1681), .ZN(n1679) );
  AOI21_X2 U2717 ( .B1(n3284), .B2(n1668), .A(n1669), .ZN(n1667) );
  NAND3_X2 U2718 ( .A1(n1658), .A2(nq[9]), .A3(n1706), .ZN(n1708) );
  AOI222_X1 U2719 ( .A1(reg_a[11]), .A2(n2416), .B1(n2352), .B2(n140), .C1(
        n2349), .C2(n3146), .ZN(n1720) );
  NAND3_X2 U2720 ( .A1(n1658), .A2(nq[5]), .A3(n1685), .ZN(n1688) );
  NAND3_X2 U2721 ( .A1(n1658), .A2(nq[7]), .A3(n1696), .ZN(n1698) );
  NOR3_X2 U2722 ( .A1(n2363), .A2(n3285), .A3(n3284), .ZN(n1669) );
  NOR3_X2 U2723 ( .A1(n2441), .A2(q[1]), .A3(n398), .ZN(n776) );
  NOR3_X2 U2724 ( .A1(n2441), .A2(q[7]), .A3(n801), .ZN(n800) );
  NOR3_X2 U2725 ( .A1(n2441), .A2(q[9]), .A3(n808), .ZN(n807) );
  NOR3_X2 U2726 ( .A1(n2441), .A2(q[5]), .A3(n794), .ZN(n793) );
  OAI21_X2 U2727 ( .B1(q[7]), .B2(n2322), .A(n802), .ZN(n804) );
  OAI21_X2 U2728 ( .B1(nq[9]), .B2(n2363), .A(n16), .ZN(n1715) );
  OAI21_X2 U2729 ( .B1(nq[5]), .B2(n2363), .A(n18), .ZN(n1695) );
  OAI21_X2 U2730 ( .B1(nq[7]), .B2(n2363), .A(n17), .ZN(n1705) );
  AND4_X2 U2731 ( .A1(n103), .A2(i_start), .A3(n968), .A4(n171), .ZN(n2332) );
  NOR3_X2 U2732 ( .A1(n1902), .A2(n1903), .A3(n1904), .ZN(n1900) );
  AOI222_X1 U2733 ( .A1(reg_b[1]), .A2(n2417), .B1(n2420), .B2(n478), .C1(
        n2413), .C2(n3120), .ZN(n774) );
  OR3_X2 U2734 ( .A1(n2417), .A2(n1976), .A3(n964), .ZN(n2333) );
  NAND3_X2 U2735 ( .A1(n645), .A2(n646), .A3(n647), .ZN(n998) );
  AOI211_X2 U2736 ( .C1(i_dividend[12]), .C2(n2426), .A(n648), .B(n633), .ZN(
        n647) );
  AOI222_X1 U2737 ( .A1(n2339), .A2(n649), .B1(n637), .B2(n650), .C1(n639), 
        .C2(n651), .ZN(n646) );
  NAND3_X2 U2738 ( .A1(n654), .A2(n655), .A3(n656), .ZN(n997) );
  AOI211_X2 U2739 ( .C1(i_dividend[13]), .C2(n2426), .A(n657), .B(n633), .ZN(
        n656) );
  AOI222_X1 U2740 ( .A1(n2339), .A2(n658), .B1(n637), .B2(n440), .C1(n639), 
        .C2(n659), .ZN(n655) );
  NAND3_X2 U2741 ( .A1(n662), .A2(n663), .A3(n664), .ZN(n996) );
  AOI211_X2 U2742 ( .C1(i_dividend[14]), .C2(n2426), .A(n665), .B(n633), .ZN(
        n664) );
  AOI222_X1 U2743 ( .A1(n2339), .A2(n669), .B1(n637), .B2(n670), .C1(n639), 
        .C2(n671), .ZN(n663) );
  NAND3_X2 U2744 ( .A1(n628), .A2(n629), .A3(n630), .ZN(n999) );
  AOI211_X2 U2745 ( .C1(i_dividend[11]), .C2(n2426), .A(n632), .B(n633), .ZN(
        n630) );
  AOI222_X1 U2746 ( .A1(n2339), .A2(n636), .B1(n637), .B2(n638), .C1(n639), 
        .C2(n640), .ZN(n629) );
  NAND3_X2 U2747 ( .A1(n1712), .A2(n1713), .A3(n1714), .ZN(n1032) );
  AOI222_X1 U2748 ( .A1(reg_a[10]), .A2(n2415), .B1(n2352), .B2(n141), .C1(
        n2349), .C2(n3144), .ZN(n1714) );
  NAND3_X2 U2749 ( .A1(n1692), .A2(n1693), .A3(n1694), .ZN(n1036) );
  AOI222_X1 U2750 ( .A1(reg_a[6]), .A2(n2417), .B1(n2353), .B2(n112), .C1(
        n2350), .C2(n3136), .ZN(n1694) );
  NAND3_X2 U2751 ( .A1(n1702), .A2(n1703), .A3(n1704), .ZN(n1034) );
  AOI222_X1 U2752 ( .A1(reg_a[8]), .A2(n2417), .B1(n2352), .B2(n143), .C1(
        n2349), .C2(n3140), .ZN(n1704) );
  NAND3_X2 U2753 ( .A1(n1682), .A2(n1683), .A3(n1684), .ZN(n1038) );
  AOI222_X1 U2754 ( .A1(reg_a[4]), .A2(n2417), .B1(n2353), .B2(n114), .C1(
        n2350), .C2(n3131), .ZN(n1684) );
  AOI222_X1 U2755 ( .A1(reg_a[31]), .A2(n2417), .B1(n2351), .B2(n119), .C1(
        n2348), .C2(n3193), .ZN(n1817) );
  NAND3_X2 U2756 ( .A1(n1658), .A2(nq[11]), .A3(n1716), .ZN(n1718) );
  BUF_X4 U2757 ( .A(i_rst), .Z(n2445) );
  BUF_X4 U2758 ( .A(i_rst), .Z(n2456) );
  BUF_X4 U2759 ( .A(i_rst), .Z(n2455) );
  BUF_X4 U2760 ( .A(i_rst), .Z(n2454) );
  BUF_X4 U2761 ( .A(i_rst), .Z(n2453) );
  BUF_X4 U2762 ( .A(i_rst), .Z(n2452) );
  BUF_X4 U2763 ( .A(i_rst), .Z(n2450) );
  BUF_X4 U2764 ( .A(i_rst), .Z(n2449) );
  BUF_X4 U2765 ( .A(i_rst), .Z(n2448) );
  BUF_X4 U2766 ( .A(i_rst), .Z(n2447) );
  BUF_X4 U2767 ( .A(i_rst), .Z(n2446) );
  BUF_X4 U2768 ( .A(i_rst), .Z(n2451) );
  BUF_X4 U2769 ( .A(i_rst), .Z(n2469) );
  BUF_X4 U2770 ( .A(i_rst), .Z(n2468) );
  BUF_X4 U2771 ( .A(i_rst), .Z(n2467) );
  BUF_X4 U2772 ( .A(i_rst), .Z(n2466) );
  BUF_X4 U2773 ( .A(i_rst), .Z(n2465) );
  BUF_X4 U2774 ( .A(i_rst), .Z(n2464) );
  BUF_X4 U2775 ( .A(i_rst), .Z(n2462) );
  BUF_X4 U2776 ( .A(i_rst), .Z(n2461) );
  BUF_X4 U2777 ( .A(i_rst), .Z(n2460) );
  BUF_X4 U2778 ( .A(i_rst), .Z(n2459) );
  BUF_X4 U2779 ( .A(i_rst), .Z(n2458) );
  BUF_X4 U2780 ( .A(i_rst), .Z(n2457) );
  BUF_X4 U2781 ( .A(i_rst), .Z(n2463) );
  AND2_X4 U2782 ( .A1(n37), .A2(n898), .ZN(n773) );
  INV_X1 U2783 ( .A(n977), .ZN(n2471) );
  NAND2_X1 U2784 ( .A1(n110), .A2(n2471), .ZN(n2470) );
endmodule

