
module s5378_bench ( blif_clk_net, blif_reset_net, n3065gat, n3066gat, 
        n3067gat, n3068gat, n3069gat, n3070gat, n3071gat, n3072gat, n3073gat, 
        n3074gat, n3075gat, n3076gat, n3077gat, n3078gat, n3079gat, n3080gat, 
        n3081gat, n3082gat, n3083gat, n3084gat, n3085gat, n3086gat, n3087gat, 
        n3088gat, n3089gat, n3090gat, n3091gat, n3092gat, n3093gat, n3094gat, 
        n3095gat, n3097gat, n3098gat, n3099gat, n3100gat, n3104gat, n3105gat, 
        n3106gat, n3107gat, n3108gat, n3109gat, n3110gat, n3111gat, n3112gat, 
        n3113gat, n3114gat, n3115gat, n3116gat, n3117gat, n3118gat, n3119gat, 
        n3120gat, n3121gat, n3122gat, n3123gat, n3124gat, n3125gat, n3126gat, 
        n3127gat, n3128gat, n3129gat, n3130gat, n3131gat, n3132gat, n3133gat, 
        n3134gat, n3135gat, n3136gat, n3137gat, n3138gat, n3139gat, n3140gat, 
        n3141gat, n3142gat, n3143gat, n3144gat, n3145gat, n3146gat, n3147gat, 
        n3148gat, n3149gat, n3150gat, n3151gat, n3152gat, test_si1, test_so1, 
        test_si2, test_so2, test_se );
  input blif_clk_net, blif_reset_net, n3065gat, n3066gat, n3067gat, n3068gat,
         n3069gat, n3070gat, n3071gat, n3072gat, n3073gat, n3074gat, n3075gat,
         n3076gat, n3077gat, n3078gat, n3079gat, n3080gat, n3081gat, n3082gat,
         n3083gat, n3084gat, n3085gat, n3086gat, n3087gat, n3088gat, n3089gat,
         n3090gat, n3091gat, n3092gat, n3093gat, n3094gat, n3095gat, n3097gat,
         n3098gat, n3099gat, n3100gat, test_si1, test_si2, test_se;
  output n3104gat, n3105gat, n3106gat, n3107gat, n3108gat, n3109gat, n3110gat,
         n3111gat, n3112gat, n3113gat, n3114gat, n3115gat, n3116gat, n3117gat,
         n3118gat, n3119gat, n3120gat, n3121gat, n3122gat, n3123gat, n3124gat,
         n3125gat, n3126gat, n3127gat, n3128gat, n3129gat, n3130gat, n3131gat,
         n3132gat, n3133gat, n3134gat, n3135gat, n3136gat, n3137gat, n3138gat,
         n3139gat, n3140gat, n3141gat, n3142gat, n3143gat, n3144gat, n3145gat,
         n3146gat, n3147gat, n3148gat, n3149gat, n3150gat, n3151gat, n3152gat,
         test_so1, test_so2;
  wire   n3140gat, n673gat, n2897gat, n398gat, n402gat, n748gat, n271gat,
         n341gat, n2472gat, n1620gat, n1827gat, n55gat, n2914gat, n2928gat,
         n2927gat, n2896gat, n2922gat, n865gat, n2894gat, n2921gat, n2895gat,
         n933gat, n834gat, n838gat, n830gat, n614gat, n504gat, n680gat,
         n2913gat, n816gat, n2920gat, n580gat, n2905gat, n824gat, n820gat,
         n2898gat, n699gat, n567gat, n2102gat, n1606gat, n1763gat, n1610gat,
         n2918gat, n2952gat, n2919gat, n2910gat, n2907gat, n931gat, n2911gat,
         n2912gat, n2909gat, n1197gat, n2908gat, n2971gat, n667gat, n2904gat,
         n2891gat, n2903gat, n2915gat, n2901gat, n2890gat, n2888gat, n2887gat,
         n2886gat, n3010gat, n3016gat, n2658gat, n2579gat, n2339gat, n2502gat,
         n2646gat, n2506gat, n2613gat, n1834gat, n1767gat, n2139gat, n1899gat,
         n2403gat, n2394gat, n2440gat, n2347gat, n1793gat, n2021gat, n1394gat,
         n1516gat, n1565gat, n2262gat, n2983gat, n1316gat, n1312gat, n1775gat,
         n1696gat, n2592gat, n1636gat, n1678gat, n2450gat, n2446gat, n2095gat,
         n2454gat, n2163gat, n2040gat, n2015gat, n2037gat, n2017gat, n2033gat,
         n463gat, n384gat, n470gat, n148gat, n1771gat, n1613gat, n1336gat,
         n1391gat, n1748gat, n1927gat, n1807gat, n1567gat, n1456gat, n1564gat,
         n1525gat, n1915gat, n1596gat, n1800gat, n1593gat, n2761gat, n2989gat,
         n2812gat, n2741gat, n2749gat, n2702gat, n2936gat, n2693gat, n2709gat,
         n2951gat, n2955gat, n2941gat, n2800gat, n2956gat, n2194gat, n2917gat,
         n2330gat, n2892gat, n2798gat, n2916gat, n2925gat, n2387gat, n2923gat,
         n2980gat, n2756gat, n2057gat, n2924gat, n2899gat, n2436gat, n2929gat,
         n2937gat, n2704gat, n2926gat, n2935gat, n1269gat, n2757gat, n2764gat,
         n2750gat, n2938gat, n2684gat, n2762gat, n2830gat, n2198gat, n1721gat,
         n2950gat, n1882gat, n2556gat, n2822gat, n2900gat, n2197gat, n2744gat,
         n1745gat, n2742gat, n2708gat, n2196gat, n2799gat, n2396gat, n1, n6,
         n7, n13, n15, n18, n19, n20, n25, n30, n31, n32, n33, n34, n37, n38,
         n39, n40, n41, n42, n46, n47, n48, n49, n50, n53, n57, n62, n63, n64,
         n65, n66, n67, n68, n69, n74, n75, n76, n79, n80, n81, n82, n83, n84,
         n85, n89, n94, n96, n97, n109, n110, n112, n113, n114, n116, n123,
         n128, n129, n132, n133, n134, n135, n136, n137, n138, n141, n142,
         n488, n489, n491, n492, n493, n494, n495, n496, n498, n499, n500,
         n502, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n5, n8, n9, n10, n11, n12, n14, n16, n17, n21, n22, n23, n24,
         n26, n27, n28, n29, n35, n36, n43, n44, n45, n51, n52, n54, n55, n56,
         n58, n59, n60, n61, n70, n71, n72, n73, n77, n78, n86, n87, n88, n90,
         n91, n92, n93, n95, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n111, n115, n117, n118, n119, n120, n121;
  assign n3152gat = 1'b1;
  assign n3115gat = 1'b1;
  assign n3112gat = 1'b1;
  assign n3139gat = n3140gat;
  assign test_so2 = n2658gat;
  assign test_so1 = n1767gat;
  assign n3123gat = n2761gat;
  assign n3105gat = n2812gat;
  assign n3117gat = n2741gat;
  assign n3119gat = n2749gat;
  assign n3113gat = n2702gat;
  assign n3131gat = n2936gat;
  assign n3114gat = n2693gat;
  assign n3111gat = n2709gat;
  assign n3129gat = n2951gat;
  assign n3130gat = n2955gat;
  assign n3137gat = n2941gat;
  assign n3143gat = n2800gat;
  assign n3133gat = n2956gat;
  assign n3108gat = n2798gat;
  assign n3142gat = n2980gat;
  assign n3141gat = n2980gat;
  assign n3121gat = n2756gat;
  assign n3134gat = n2937gat;
  assign n3151gat = n2704gat;
  assign n3135gat = n2935gat;
  assign n3116gat = n1269gat;
  assign n3122gat = n2757gat;
  assign n3125gat = n2764gat;
  assign n3120gat = n2750gat;
  assign n3132gat = n2938gat;
  assign n3150gat = n2684gat;
  assign n3124gat = n2762gat;
  assign n3147gat = n2830gat;
  assign n3138gat = n1721gat;
  assign n3136gat = n2950gat;
  assign n3104gat = n2822gat;
  assign n3144gat = n2744gat;
  assign n3107gat = n1745gat;
  assign n3118gat = n2742gat;
  assign n3110gat = n2708gat;
  assign n3109gat = n2799gat;

  INV_X4 U535 ( .A(blif_reset_net), .ZN(n559) );
  INV_X4 U536 ( .A(blif_reset_net), .ZN(n564) );
  INV_X4 U537 ( .A(n573), .ZN(n565) );
  INV_X4 U538 ( .A(n574), .ZN(n566) );
  INV_X4 U539 ( .A(blif_reset_net), .ZN(n561) );
  INV_X4 U540 ( .A(n573), .ZN(n563) );
  INV_X4 U541 ( .A(n574), .ZN(n562) );
  INV_X4 U542 ( .A(blif_reset_net), .ZN(n560) );
  INV_X4 U543 ( .A(n574), .ZN(n569) );
  INV_X4 U544 ( .A(n573), .ZN(n570) );
  INV_X4 U545 ( .A(n574), .ZN(n568) );
  INV_X4 U546 ( .A(n573), .ZN(n571) );
  INV_X4 U547 ( .A(n574), .ZN(n567) );
  INV_X4 U548 ( .A(n573), .ZN(n572) );
  INV_X4 U549 ( .A(n1), .ZN(n573) );
  INV_X4 U550 ( .A(n1), .ZN(n574) );
  INV_X1 U551 ( .A(n575), .ZN(n94) );
  INV_X1 U552 ( .A(n576), .ZN(n7) );
  OAI211_X1 U553 ( .C1(n116), .C2(n1312gat), .A(n2017gat), .B(n577), .ZN(n576)
         );
  MUX2_X1 U554 ( .A(n578), .B(n579), .S(n580), .Z(n502) );
  NOR3_X1 U555 ( .A1(n581), .A2(n582), .A3(n583), .ZN(n579) );
  NAND3_X1 U556 ( .A1(n3087gat), .A2(n510), .A3(n584), .ZN(n581) );
  AND3_X1 U557 ( .A1(n3094gat), .A2(n585), .A3(n586), .ZN(n578) );
  NOR3_X1 U558 ( .A1(n587), .A2(n532), .A3(n588), .ZN(n499) );
  NAND2_X1 U559 ( .A1(n18), .A2(n589), .ZN(n495) );
  XOR2_X1 U560 ( .A(n963), .B(n590), .Z(n589) );
  AND3_X1 U561 ( .A1(n591), .A2(n532), .A3(n587), .ZN(n590) );
  NAND2_X1 U562 ( .A1(n19), .A2(n592), .ZN(n494) );
  XOR2_X1 U563 ( .A(n962), .B(n593), .Z(n592) );
  AOI211_X1 U564 ( .C1(n2403gat), .C2(n505), .A(n2440gat), .B(n594), .ZN(n593)
         );
  NAND2_X1 U565 ( .A1(n20), .A2(n595), .ZN(n493) );
  XOR2_X1 U566 ( .A(n961), .B(n596), .Z(n595) );
  NOR2_X1 U567 ( .A1(n2262gat), .A2(n997), .ZN(n596) );
  NAND3_X1 U568 ( .A1(n597), .A2(n598), .A3(n599), .ZN(n488) );
  NOR4_X1 U569 ( .A1(n600), .A2(n136), .A3(n545), .A4(n129), .ZN(n3146gat) );
  NAND4_X1 U570 ( .A1(n2033gat), .A2(n2095gat), .A3(n2037gat), .A4(n601), .ZN(
        n600) );
  NAND3_X1 U571 ( .A1(n510), .A2(n549), .A3(n602), .ZN(n601) );
  AOI21_X1 U572 ( .B1(n602), .B2(n549), .A(n6), .ZN(n3145gat) );
  INV_X1 U573 ( .A(n598), .ZN(n6) );
  NOR2_X1 U574 ( .A1(n489), .A2(n492), .ZN(n598) );
  INV_X1 U575 ( .A(n603), .ZN(n492) );
  NAND2_X1 U576 ( .A1(n604), .A2(n605), .ZN(n489) );
  NAND2_X1 U577 ( .A1(n606), .A2(n607), .ZN(n3140gat) );
  OAI211_X1 U578 ( .C1(n608), .C2(n32), .A(n116), .B(n609), .ZN(n607) );
  NOR2_X1 U579 ( .A1(n3106gat), .A2(n3098gat), .ZN(n609) );
  AND3_X1 U580 ( .A1(n610), .A2(n546), .A3(n3097gat), .ZN(n608) );
  MUX2_X1 U581 ( .A(n611), .B(n612), .S(n2989gat), .Z(n606) );
  INV_X1 U582 ( .A(n613), .ZN(n612) );
  OAI22_X1 U583 ( .A1(n614), .A2(n982), .B1(n1678gat), .B2(n1008), .ZN(n613)
         );
  INV_X1 U584 ( .A(n615), .ZN(n614) );
  OAI33_X1 U585 ( .A1(n555), .A2(n616), .A3(n109), .B1(n521), .B2(n617), .B3(
        n618), .ZN(n615) );
  NOR2_X1 U586 ( .A1(n619), .A2(n620), .ZN(n611) );
  MUX2_X1 U587 ( .A(n621), .B(n960), .S(n1596gat), .Z(n620) );
  AOI21_X1 U588 ( .B1(n604), .B2(n109), .A(n1678gat), .ZN(n621) );
  NOR3_X1 U589 ( .A1(n1525gat), .A2(n1394gat), .A3(n622), .ZN(n619) );
  NAND2_X1 U590 ( .A1(n623), .A2(n624), .ZN(n3016gat) );
  NOR4_X1 U591 ( .A1(n964), .A2(n965), .A3(n966), .A4(n967), .ZN(n624) );
  NOR4_X1 U592 ( .A1(n968), .A2(n969), .A3(n970), .A4(n3090gat), .ZN(n623) );
  NOR3_X1 U593 ( .A1(n625), .A2(n626), .A3(n627), .ZN(n2983gat) );
  AOI21_X1 U594 ( .B1(n972), .B2(n628), .A(n971), .ZN(n627) );
  MUX2_X1 U595 ( .A(n629), .B(n630), .S(n2989gat), .Z(n2980gat) );
  OAI22_X1 U596 ( .A1(n142), .A2(n1807gat), .B1(n631), .B2(n1456gat), .ZN(n630) );
  AOI21_X1 U597 ( .B1(n142), .B2(n632), .A(n3149gat), .ZN(n631) );
  INV_X1 U598 ( .A(n618), .ZN(n632) );
  NOR2_X1 U599 ( .A1(n633), .A2(n491), .ZN(n618) );
  OAI21_X1 U600 ( .B1(n634), .B2(n1748gat), .A(n635), .ZN(n629) );
  NAND3_X1 U601 ( .A1(n491), .A2(n109), .A3(n973), .ZN(n635) );
  AOI211_X1 U602 ( .C1(n491), .C2(n1336gat), .A(n633), .B(n3149gat), .ZN(n634)
         );
  OAI22_X1 U603 ( .A1(n636), .A2(n637), .B1(n638), .B2(n639), .ZN(n2956gat) );
  AOI222_X1 U604 ( .A1(n640), .A2(n42), .B1(n641), .B2(n519), .C1(n642), .C2(
        n551), .ZN(n639) );
  OAI22_X1 U605 ( .A1(n637), .A2(n643), .B1(n638), .B2(n644), .ZN(n2955gat) );
  AOI222_X1 U606 ( .A1(n640), .A2(n38), .B1(n641), .B2(n517), .C1(n642), .C2(
        n75), .ZN(n644) );
  OAI21_X1 U607 ( .B1(n645), .B2(n646), .A(n647), .ZN(n2952gat) );
  OAI22_X1 U608 ( .A1(n638), .A2(n648), .B1(n637), .B2(n649), .ZN(n2951gat) );
  AOI222_X1 U609 ( .A1(n640), .A2(n41), .B1(n641), .B2(n516), .C1(n642), .C2(
        n1269gat), .ZN(n648) );
  OAI222_X1 U610 ( .A1(n637), .A2(n650), .B1(n531), .B2(n651), .C1(n504), .C2(
        n652), .ZN(n2950gat) );
  OAI222_X1 U611 ( .A1(n637), .A2(n653), .B1(n556), .B2(n651), .C1(n511), .C2(
        n652), .ZN(n2941gat) );
  OAI22_X1 U612 ( .A1(n637), .A2(n654), .B1(n638), .B2(n655), .ZN(n2938gat) );
  AOI222_X1 U613 ( .A1(n640), .A2(n39), .B1(n641), .B2(n25), .C1(n642), .C2(
        n76), .ZN(n655) );
  OAI222_X1 U614 ( .A1(n637), .A2(n656), .B1(n539), .B2(n651), .C1(n398gat), 
        .C2(n652), .ZN(n2937gat) );
  OAI22_X1 U615 ( .A1(n637), .A2(n657), .B1(n638), .B2(n658), .ZN(n2936gat) );
  AOI222_X1 U616 ( .A1(n640), .A2(n40), .B1(n641), .B2(n991), .C1(n642), .C2(
        n1005), .ZN(n658) );
  INV_X1 U617 ( .A(n659), .ZN(n638) );
  OAI222_X1 U618 ( .A1(n637), .A2(n660), .B1(n530), .B2(n651), .C1(n402gat), 
        .C2(n652), .ZN(n2935gat) );
  OAI21_X1 U619 ( .B1(n640), .B2(n641), .A(n659), .ZN(n652) );
  NAND2_X1 U620 ( .A1(n642), .A2(n659), .ZN(n651) );
  OAI21_X1 U621 ( .B1(n580), .B2(n661), .A(n662), .ZN(n659) );
  INV_X1 U622 ( .A(n663), .ZN(n637) );
  OAI21_X1 U623 ( .B1(n3088gat), .B2(n661), .A(n664), .ZN(n663) );
  NAND3_X1 U624 ( .A1(n665), .A2(n3086gat), .A3(n666), .ZN(n664) );
  OAI21_X1 U625 ( .B1(n667), .B2(n668), .A(n584), .ZN(n661) );
  OAI222_X1 U626 ( .A1(n669), .A2(n670), .B1(n671), .B2(n672), .C1(n673), .C2(
        n674), .ZN(n2929gat) );
  INV_X1 U627 ( .A(n3081gat), .ZN(n674) );
  XNOR2_X1 U628 ( .A(n675), .B(n978), .ZN(n671) );
  INV_X1 U629 ( .A(n676), .ZN(n2928gat) );
  INV_X1 U630 ( .A(n677), .ZN(n2927gat) );
  MUX2_X1 U631 ( .A(n3073gat), .B(n678), .S(n679), .Z(n2926gat) );
  XOR2_X1 U632 ( .A(n470gat), .B(n680), .Z(n678) );
  NAND2_X1 U633 ( .A1(n681), .A2(n682), .ZN(n680) );
  OAI21_X1 U634 ( .B1(n974), .B2(n975), .A(n979), .ZN(n682) );
  OAI222_X1 U635 ( .A1(n669), .A2(n683), .B1(n684), .B2(n672), .C1(n673), .C2(
        n685), .ZN(n2925gat) );
  INV_X1 U636 ( .A(n3082gat), .ZN(n685) );
  XOR2_X1 U637 ( .A(n463gat), .B(n686), .Z(n684) );
  AND2_X1 U638 ( .A1(n687), .A2(n675), .ZN(n686) );
  OAI21_X1 U639 ( .B1(n977), .B2(n976), .A(n978), .ZN(n687) );
  MUX2_X1 U640 ( .A(n3066gat), .B(n688), .S(n679), .Z(n2924gat) );
  XOR2_X1 U641 ( .A(n974), .B(n689), .Z(n688) );
  MUX2_X1 U642 ( .A(n3065gat), .B(n690), .S(n679), .Z(n2923gat) );
  XOR2_X1 U643 ( .A(n148gat), .B(n691), .Z(n690) );
  NAND2_X1 U644 ( .A1(n689), .A2(n974), .ZN(n691) );
  NOR2_X1 U645 ( .A1(n692), .A2(n975), .ZN(n689) );
  INV_X1 U646 ( .A(n693), .ZN(n2922gat) );
  INV_X1 U647 ( .A(n694), .ZN(n2921gat) );
  OAI22_X1 U648 ( .A1(n673), .A2(n695), .B1(n646), .B2(n669), .ZN(n2920gat) );
  INV_X1 U649 ( .A(n3067gat), .ZN(n646) );
  INV_X1 U650 ( .A(n3076gat), .ZN(n695) );
  OAI21_X1 U651 ( .B1(n645), .B2(n696), .A(n647), .ZN(n2919gat) );
  OAI21_X1 U652 ( .B1(n645), .B2(n697), .A(n647), .ZN(n2918gat) );
  MUX2_X1 U653 ( .A(n3067gat), .B(n698), .S(n679), .Z(n2917gat) );
  XOR2_X1 U654 ( .A(n692), .B(n975), .Z(n698) );
  NAND2_X1 U655 ( .A1(n681), .A2(n979), .ZN(n692) );
  OAI222_X1 U656 ( .A1(n669), .A2(n699), .B1(n700), .B2(n672), .C1(n673), .C2(
        n701), .ZN(n2916gat) );
  INV_X1 U657 ( .A(n3079gat), .ZN(n701) );
  XNOR2_X1 U658 ( .A(n702), .B(n536), .ZN(n700) );
  NAND2_X1 U659 ( .A1(n647), .A2(n677), .ZN(n2915gat) );
  AOI22_X1 U660 ( .A1(n3095gat), .A2(n3075gat), .B1(n3093gat), .B2(n3066gat), 
        .ZN(n677) );
  INV_X1 U661 ( .A(n703), .ZN(n2914gat) );
  OAI22_X1 U662 ( .A1(n673), .A2(n704), .B1(n669), .B2(n697), .ZN(n2913gat) );
  INV_X1 U663 ( .A(n3065gat), .ZN(n697) );
  INV_X1 U664 ( .A(n3074gat), .ZN(n704) );
  OAI21_X1 U665 ( .B1(n645), .B2(n699), .A(n647), .ZN(n2912gat) );
  INV_X1 U666 ( .A(n3070gat), .ZN(n699) );
  OAI21_X1 U667 ( .B1(n645), .B2(n705), .A(n647), .ZN(n2911gat) );
  OAI21_X1 U668 ( .B1(n645), .B2(n706), .A(n647), .ZN(n2910gat) );
  OAI21_X1 U669 ( .B1(n645), .B2(n707), .A(n647), .ZN(n2909gat) );
  OAI21_X1 U670 ( .B1(n645), .B2(n683), .A(n647), .ZN(n2908gat) );
  INV_X1 U671 ( .A(n3073gat), .ZN(n683) );
  OAI21_X1 U672 ( .B1(n645), .B2(n670), .A(n647), .ZN(n2907gat) );
  INV_X1 U673 ( .A(n3072gat), .ZN(n670) );
  INV_X1 U674 ( .A(n708), .ZN(n645) );
  OAI33_X1 U675 ( .A1(n709), .A2(n710), .A3(n582), .B1(n711), .B2(n712), .B3(
        n713), .ZN(n708) );
  OAI22_X1 U676 ( .A1(n673), .A2(n714), .B1(n669), .B2(n696), .ZN(n2905gat) );
  INV_X1 U677 ( .A(n3066gat), .ZN(n696) );
  INV_X1 U678 ( .A(n3075gat), .ZN(n714) );
  NAND2_X1 U679 ( .A1(n647), .A2(n693), .ZN(n2904gat) );
  AOI22_X1 U680 ( .A1(n3095gat), .A2(n3082gat), .B1(n3093gat), .B2(n3073gat), 
        .ZN(n693) );
  NAND2_X1 U681 ( .A1(n647), .A2(n676), .ZN(n2903gat) );
  AOI22_X1 U682 ( .A1(n3095gat), .A2(n3076gat), .B1(n3093gat), .B2(n3067gat), 
        .ZN(n676) );
  NAND2_X1 U683 ( .A1(n647), .A2(n715), .ZN(n2901gat) );
  OAI222_X1 U684 ( .A1(n669), .A2(n706), .B1(n672), .B2(n716), .C1(n673), .C2(
        n717), .ZN(n2900gat) );
  INV_X1 U685 ( .A(n3080gat), .ZN(n717) );
  XNOR2_X1 U686 ( .A(n542), .B(n718), .ZN(n716) );
  INV_X1 U687 ( .A(n3071gat), .ZN(n706) );
  OAI222_X1 U688 ( .A1(n669), .A2(n707), .B1(n719), .B2(n672), .C1(n673), .C2(
        n720), .ZN(n2899gat) );
  INV_X1 U689 ( .A(n3078gat), .ZN(n720) );
  NAND2_X1 U690 ( .A1(n673), .A2(n669), .ZN(n672) );
  XOR2_X1 U691 ( .A(n384gat), .B(n721), .Z(n719) );
  NOR2_X1 U692 ( .A1(n536), .A2(n702), .ZN(n721) );
  NAND2_X1 U693 ( .A1(n718), .A2(n542), .ZN(n702) );
  AND2_X1 U694 ( .A1(n675), .A2(n978), .ZN(n718) );
  INV_X1 U695 ( .A(n3069gat), .ZN(n707) );
  OAI22_X1 U696 ( .A1(n673), .A2(n722), .B1(n669), .B2(n705), .ZN(n2898gat) );
  INV_X1 U697 ( .A(n3068gat), .ZN(n705) );
  NAND3_X1 U698 ( .A1(n723), .A2(n724), .A3(n725), .ZN(n669) );
  NOR3_X1 U699 ( .A1(n726), .A2(n3088gat), .A3(n3086gat), .ZN(n725) );
  INV_X1 U700 ( .A(n3077gat), .ZN(n722) );
  INV_X1 U701 ( .A(n727), .ZN(n2897gat) );
  INV_X1 U702 ( .A(n715), .ZN(n2896gat) );
  AOI22_X1 U703 ( .A1(n3095gat), .A2(n3080gat), .B1(n3093gat), .B2(n3071gat), 
        .ZN(n715) );
  INV_X1 U704 ( .A(n728), .ZN(n2895gat) );
  INV_X1 U705 ( .A(n729), .ZN(n2894gat) );
  MUX2_X1 U706 ( .A(n3068gat), .B(n730), .S(n679), .Z(n2892gat) );
  AND2_X1 U707 ( .A1(n673), .A2(n731), .ZN(n679) );
  NAND4_X1 U708 ( .A1(n723), .A2(n666), .A3(n724), .A4(n710), .ZN(n731) );
  NAND4_X1 U709 ( .A1(n3094gat), .A2(n586), .A3(n3088gat), .A4(n712), .ZN(n673) );
  XOR2_X1 U710 ( .A(n979), .B(n681), .Z(n730) );
  NAND2_X1 U711 ( .A1(n647), .A2(n703), .ZN(n2891gat) );
  AOI22_X1 U712 ( .A1(n3095gat), .A2(n3074gat), .B1(n3093gat), .B2(n3065gat), 
        .ZN(n703) );
  NAND2_X1 U713 ( .A1(n647), .A2(n727), .ZN(n2890gat) );
  AOI22_X1 U714 ( .A1(n3095gat), .A2(n3081gat), .B1(n3093gat), .B2(n3072gat), 
        .ZN(n727) );
  NAND2_X1 U715 ( .A1(n647), .A2(n729), .ZN(n2888gat) );
  AOI22_X1 U716 ( .A1(n3095gat), .A2(n3077gat), .B1(n3093gat), .B2(n3068gat), 
        .ZN(n729) );
  NAND2_X1 U717 ( .A1(n647), .A2(n694), .ZN(n2887gat) );
  AOI22_X1 U718 ( .A1(n3095gat), .A2(n3079gat), .B1(n3093gat), .B2(n3070gat), 
        .ZN(n694) );
  NAND2_X1 U719 ( .A1(n647), .A2(n728), .ZN(n2886gat) );
  AOI22_X1 U720 ( .A1(n3095gat), .A2(n3078gat), .B1(n3093gat), .B2(n3069gat), 
        .ZN(n728) );
  NAND4_X1 U721 ( .A1(n732), .A2(n538), .A3(n733), .A4(n734), .ZN(n647) );
  AND4_X1 U722 ( .A1(n64), .A2(n67), .A3(n735), .A4(n736), .ZN(n734) );
  INV_X1 U723 ( .A(n737), .ZN(n736) );
  MUX2_X1 U724 ( .A(n527), .B(n74), .S(n512), .Z(n737) );
  MUX2_X1 U725 ( .A(n74), .B(n527), .S(n65), .Z(n735) );
  AOI21_X1 U726 ( .B1(n738), .B2(n62), .A(n622), .ZN(n733) );
  INV_X1 U727 ( .A(n491), .ZN(n622) );
  NAND2_X1 U728 ( .A1(n605), .A2(n603), .ZN(n491) );
  AND2_X1 U729 ( .A1(n739), .A2(n740), .ZN(n605) );
  NAND4_X1 U730 ( .A1(n402gat), .A2(n741), .A3(n543), .A4(n504), .ZN(n740) );
  INV_X1 U731 ( .A(n617), .ZN(n732) );
  NOR4_X1 U732 ( .A1(n534), .A2(n508), .A3(n742), .A4(n53), .ZN(n617) );
  OAI211_X1 U733 ( .C1(n743), .C2(n744), .A(n745), .B(n746), .ZN(n2822gat) );
  OR3_X1 U734 ( .A1(n712), .A2(n586), .A3(n711), .ZN(n745) );
  INV_X1 U735 ( .A(n713), .ZN(n586) );
  OR2_X1 U736 ( .A1(n747), .A2(n748), .ZN(n2812gat) );
  OAI33_X1 U737 ( .A1(n709), .A2(n3086gat), .A3(n582), .B1(n711), .B2(n585), 
        .B3(n713), .ZN(n748) );
  NAND2_X1 U738 ( .A1(n3094gat), .A2(n580), .ZN(n711) );
  INV_X1 U739 ( .A(n724), .ZN(n582) );
  NOR2_X1 U740 ( .A1(n749), .A2(n743), .ZN(n724) );
  NOR2_X1 U741 ( .A1(n3091gat), .A2(n3092gat), .ZN(n743) );
  NAND2_X1 U742 ( .A1(n750), .A2(n2613gat), .ZN(n2800gat) );
  NAND2_X1 U743 ( .A1(n554), .A2(n751), .ZN(n2799gat) );
  NAND2_X1 U744 ( .A1(n752), .A2(n558), .ZN(n2798gat) );
  OAI21_X1 U745 ( .B1(n649), .B2(n662), .A(n2646gat), .ZN(n2764gat) );
  AOI221_X1 U746 ( .B1(n980), .B2(n641), .C1(n47), .C2(n640), .A(n753), .ZN(
        n649) );
  INV_X1 U747 ( .A(n754), .ZN(n753) );
  AOI222_X1 U748 ( .A1(n755), .A2(n516), .B1(n756), .B2(n757), .C1(n642), .C2(
        n758), .ZN(n754) );
  AOI21_X1 U749 ( .B1(n759), .B2(n525), .A(n760), .ZN(n756) );
  OAI21_X1 U750 ( .B1(n653), .B2(n662), .A(n2971gat), .ZN(n2762gat) );
  XNOR2_X1 U751 ( .A(n1197gat), .B(n1269gat), .ZN(n2971gat) );
  AOI221_X1 U752 ( .B1(n1007), .B2(n755), .C1(n989), .C2(n642), .A(n761), .ZN(
        n653) );
  INV_X1 U753 ( .A(n762), .ZN(n761) );
  AOI22_X1 U754 ( .A1(n763), .A2(n525), .B1(n640), .B2(n48), .ZN(n762) );
  OAI21_X1 U755 ( .B1(n650), .B2(n662), .A(n3010gat), .ZN(n2761gat) );
  XNOR2_X1 U756 ( .A(n667gat), .B(n758), .ZN(n3010gat) );
  AOI221_X1 U757 ( .B1(n1006), .B2(n755), .C1(n985), .C2(n641), .A(n764), .ZN(
        n650) );
  INV_X1 U758 ( .A(n765), .ZN(n764) );
  AOI22_X1 U759 ( .A1(n642), .A2(n81), .B1(n640), .B2(n46), .ZN(n765) );
  OAI21_X1 U760 ( .B1(n660), .B2(n662), .A(n504gat), .ZN(n2757gat) );
  XOR2_X1 U761 ( .A(n766), .B(n767), .Z(n504gat) );
  XOR2_X1 U762 ( .A(n768), .B(n769), .Z(n767) );
  XNOR2_X1 U763 ( .A(n39), .B(n770), .ZN(n769) );
  MUX2_X1 U764 ( .A(n771), .B(n772), .S(n42), .Z(n768) );
  XNOR2_X1 U765 ( .A(n830gat), .B(n773), .ZN(n766) );
  XNOR2_X1 U766 ( .A(n40), .B(n834gat), .ZN(n773) );
  AOI221_X1 U767 ( .B1(n507), .B2(n755), .C1(n37), .C2(n641), .A(n774), .ZN(
        n660) );
  INV_X1 U768 ( .A(n775), .ZN(n774) );
  AOI22_X1 U769 ( .A1(n642), .A2(n82), .B1(n640), .B2(n49), .ZN(n775) );
  OAI21_X1 U770 ( .B1(n656), .B2(n662), .A(n567gat), .ZN(n2756gat) );
  XNOR2_X1 U771 ( .A(n816gat), .B(n776), .ZN(n567gat) );
  XOR2_X1 U772 ( .A(n777), .B(n778), .Z(n776) );
  XOR2_X1 U773 ( .A(n779), .B(n780), .Z(n778) );
  XNOR2_X1 U774 ( .A(n540), .B(n580gat), .ZN(n780) );
  XNOR2_X1 U775 ( .A(n820gat), .B(n50), .ZN(n779) );
  XOR2_X1 U776 ( .A(n781), .B(n782), .Z(n777) );
  XNOR2_X1 U777 ( .A(n48), .B(n824gat), .ZN(n782) );
  XNOR2_X1 U778 ( .A(n49), .B(n984), .ZN(n781) );
  AOI221_X1 U779 ( .B1(n523), .B2(n755), .C1(n983), .C2(n641), .A(n783), .ZN(
        n656) );
  INV_X1 U780 ( .A(n784), .ZN(n783) );
  AOI22_X1 U781 ( .A1(n642), .A2(n83), .B1(n640), .B2(n50), .ZN(n784) );
  OAI21_X1 U782 ( .B1(n636), .B2(n662), .A(n55gat), .ZN(n2750gat) );
  INV_X1 U783 ( .A(n785), .ZN(n636) );
  OAI221_X1 U784 ( .B1(n341gat), .B2(n786), .C1(n865gat), .C2(n787), .A(n788), 
        .ZN(n785) );
  AOI22_X1 U785 ( .A1(n642), .A2(n987), .B1(n640), .B2(n984), .ZN(n788) );
  OAI21_X1 U786 ( .B1(n654), .B2(n662), .A(n933gat), .ZN(n2749gat) );
  XNOR2_X1 U787 ( .A(n537), .B(n789), .ZN(n933gat) );
  XOR2_X1 U788 ( .A(n790), .B(n791), .Z(n789) );
  XOR2_X1 U789 ( .A(n792), .B(n793), .Z(n791) );
  XOR2_X1 U790 ( .A(n37), .B(n34), .Z(n793) );
  XNOR2_X1 U791 ( .A(n865gat), .B(n525), .ZN(n792) );
  XOR2_X1 U792 ( .A(n794), .B(n795), .Z(n790) );
  XNOR2_X1 U793 ( .A(n985), .B(n515), .ZN(n795) );
  XNOR2_X1 U794 ( .A(n980), .B(n535), .ZN(n794) );
  AOI221_X1 U795 ( .B1(n25), .B2(n755), .C1(n515), .C2(n641), .A(n796), .ZN(
        n654) );
  INV_X1 U796 ( .A(n797), .ZN(n796) );
  AOI22_X1 U797 ( .A1(n642), .A2(n988), .B1(n640), .B2(n547), .ZN(n797) );
  NAND2_X1 U798 ( .A1(n750), .A2(n2579gat), .ZN(n2744gat) );
  NOR3_X1 U799 ( .A1(n798), .A2(n799), .A3(n800), .ZN(n750) );
  OAI33_X1 U800 ( .A1(n801), .A2(n1394gat), .A3(n616), .B1(n802), .B2(n604), 
        .B3(n534), .ZN(n800) );
  INV_X1 U801 ( .A(n633), .ZN(n604) );
  MUX2_X1 U802 ( .A(n803), .B(n804), .S(n508), .Z(n802) );
  AOI221_X1 U803 ( .B1(n53), .B2(n805), .C1(n806), .C2(n57), .A(n807), .ZN(
        n804) );
  INV_X1 U804 ( .A(n808), .ZN(n807) );
  AOI22_X1 U805 ( .A1(n79), .A2(n809), .B1(n80), .B2(n738), .ZN(n808) );
  MUX2_X1 U806 ( .A(n810), .B(n811), .S(n506), .Z(n806) );
  MUX2_X1 U807 ( .A(n988), .B(n81), .S(n53), .Z(n811) );
  MUX2_X1 U808 ( .A(n987), .B(n989), .S(n53), .Z(n810) );
  OAI22_X1 U809 ( .A1(n520), .A2(n812), .B1(n541), .B2(n813), .ZN(n805) );
  NAND2_X1 U810 ( .A1(n814), .A2(n809), .ZN(n803) );
  XNOR2_X1 U811 ( .A(n815), .B(n758), .ZN(n814) );
  XOR2_X1 U812 ( .A(n816), .B(n817), .Z(n758) );
  XOR2_X1 U813 ( .A(n818), .B(n819), .Z(n817) );
  XNOR2_X1 U814 ( .A(n989), .B(n520), .ZN(n819) );
  XOR2_X1 U815 ( .A(n987), .B(n988), .Z(n818) );
  XOR2_X1 U816 ( .A(n820), .B(n821), .Z(n816) );
  XNOR2_X1 U817 ( .A(n541), .B(n81), .ZN(n821) );
  XNOR2_X1 U818 ( .A(n79), .B(n80), .ZN(n820) );
  MUX2_X1 U819 ( .A(n1678gat), .B(n982), .S(n2989gat), .Z(n801) );
  NOR2_X1 U820 ( .A1(n981), .A2(n822), .ZN(n799) );
  AOI21_X1 U821 ( .B1(n823), .B2(n824), .A(n825), .ZN(n822) );
  AOI211_X1 U822 ( .C1(n826), .C2(n827), .A(n508), .B(n64), .ZN(n825) );
  MUX2_X1 U823 ( .A(n828), .B(n829), .S(n3149gat), .Z(n827) );
  AOI22_X1 U824 ( .A1(n738), .A2(n525), .B1(n809), .B2(n985), .ZN(n829) );
  AOI22_X1 U825 ( .A1(n738), .A2(n48), .B1(n809), .B2(n46), .ZN(n828) );
  MUX2_X1 U826 ( .A(n830), .B(n831), .S(n53), .Z(n826) );
  OAI221_X1 U827 ( .B1(n39), .B2(n832), .C1(n25), .C2(n833), .A(n834), .ZN(
        n831) );
  AOI221_X1 U828 ( .B1(n835), .B2(n614gat), .C1(n836), .C2(n341gat), .A(n57), 
        .ZN(n834) );
  OAI211_X1 U829 ( .C1(n517), .C2(n833), .A(n57), .B(n837), .ZN(n830) );
  AOI222_X1 U830 ( .A1(n838), .A2(n834gat), .B1(n836), .B2(n544), .C1(n835), 
        .C2(n838gat), .ZN(n837) );
  NAND3_X1 U831 ( .A1(n839), .A2(n840), .A3(n841), .ZN(n824) );
  MUX2_X1 U832 ( .A(n842), .B(n843), .S(n53), .Z(n841) );
  MUX2_X1 U833 ( .A(n844), .B(n845), .S(n524), .Z(n843) );
  OAI221_X1 U834 ( .B1(n547), .B2(n832), .C1(n515), .C2(n833), .A(n846), .ZN(
        n845) );
  AOI22_X1 U835 ( .A1(n836), .A2(n865gat), .B1(n835), .B2(n553), .ZN(n846) );
  AOI221_X1 U836 ( .B1(n836), .B2(n37), .C1(n835), .C2(n49), .A(n847), .ZN(
        n844) );
  OAI22_X1 U837 ( .A1(n535), .A2(n833), .B1(n699gat), .B2(n832), .ZN(n847) );
  INV_X1 U838 ( .A(n838), .ZN(n832) );
  OAI211_X1 U839 ( .C1(n34), .C2(n833), .A(n57), .B(n848), .ZN(n842) );
  AOI222_X1 U840 ( .A1(n838), .A2(n680gat), .B1(n836), .B2(n537), .C1(n835), 
        .C2(n580gat), .ZN(n848) );
  NOR2_X1 U841 ( .A1(n506), .A2(n3149gat), .ZN(n835) );
  NOR2_X1 U842 ( .A1(n506), .A2(n616), .ZN(n836) );
  INV_X1 U843 ( .A(n3149gat), .ZN(n616) );
  NOR2_X1 U844 ( .A1(n3149gat), .A2(n63), .ZN(n838) );
  NAND2_X1 U845 ( .A1(n506), .A2(n3149gat), .ZN(n833) );
  OAI21_X1 U846 ( .B1(n849), .B2(n633), .A(n738), .ZN(n840) );
  NAND2_X1 U847 ( .A1(n815), .A2(n850), .ZN(n633) );
  NAND3_X1 U848 ( .A1(n851), .A2(n852), .A3(n402gat), .ZN(n850) );
  NAND2_X1 U849 ( .A1(n853), .A2(n402gat), .ZN(n815) );
  OAI21_X1 U850 ( .B1(n849), .B2(n986), .A(n809), .ZN(n839) );
  INV_X1 U851 ( .A(n739), .ZN(n849) );
  NAND4_X1 U852 ( .A1(n402gat), .A2(n851), .A3(n523), .A4(n504), .ZN(n739) );
  NOR3_X1 U853 ( .A1(n2592gat), .A2(n673gat), .A3(n3106gat), .ZN(n798) );
  OAI21_X1 U854 ( .B1(n657), .B2(n662), .A(n55gat), .ZN(n2742gat) );
  XOR2_X1 U855 ( .A(n854), .B(n855), .Z(n55gat) );
  XOR2_X1 U856 ( .A(n856), .B(n857), .Z(n855) );
  XOR2_X1 U857 ( .A(n25), .B(n770), .Z(n857) );
  XNOR2_X1 U858 ( .A(n511), .B(n1006), .ZN(n770) );
  MUX2_X1 U859 ( .A(n771), .B(n772), .S(n519), .Z(n856) );
  XNOR2_X1 U860 ( .A(n398gat), .B(n402gat), .ZN(n772) );
  OAI21_X1 U861 ( .B1(n398gat), .B2(n507), .A(n858), .ZN(n771) );
  XNOR2_X1 U862 ( .A(n271gat), .B(n859), .ZN(n854) );
  XNOR2_X1 U863 ( .A(n516), .B(n991), .ZN(n859) );
  AOI221_X1 U864 ( .B1(n991), .B2(n755), .C1(n990), .C2(n641), .A(n860), .ZN(
        n657) );
  INV_X1 U865 ( .A(n861), .ZN(n860) );
  AOI22_X1 U866 ( .A1(n642), .A2(n80), .B1(n640), .B2(n552), .ZN(n861) );
  OAI21_X1 U867 ( .B1(n643), .B2(n662), .A(n748gat), .ZN(n2741gat) );
  XNOR2_X1 U868 ( .A(n862), .B(n863), .ZN(n748gat) );
  MUX2_X1 U869 ( .A(n864), .B(n865), .S(n3089gat), .Z(n863) );
  XNOR2_X1 U870 ( .A(n580), .B(n3087gat), .ZN(n865) );
  OAI21_X1 U871 ( .B1(n3088gat), .B2(n3087gat), .A(n866), .ZN(n864) );
  INV_X1 U872 ( .A(n666), .ZN(n866) );
  NOR2_X1 U873 ( .A1(n726), .A2(n580), .ZN(n666) );
  XNOR2_X1 U874 ( .A(n867), .B(n710), .ZN(n862) );
  MUX2_X1 U875 ( .A(n868), .B(n869), .S(n749), .Z(n867) );
  XNOR2_X1 U876 ( .A(n3083gat), .B(n3084gat), .ZN(n869) );
  AOI21_X1 U877 ( .B1(n3083gat), .B2(n3084gat), .A(n584), .ZN(n868) );
  OAI21_X1 U878 ( .B1(n3087gat), .B2(n3086gat), .A(n665), .ZN(n662) );
  AOI221_X1 U879 ( .B1(n517), .B2(n755), .C1(n34), .C2(n641), .A(n870), .ZN(
        n643) );
  INV_X1 U880 ( .A(n871), .ZN(n870) );
  AOI22_X1 U881 ( .A1(n642), .A2(n79), .B1(n640), .B2(n540), .ZN(n871) );
  NOR2_X1 U882 ( .A1(n759), .A2(n757), .ZN(n640) );
  INV_X1 U883 ( .A(n872), .ZN(n759) );
  AND2_X1 U884 ( .A1(n757), .A2(n760), .ZN(n642) );
  INV_X1 U885 ( .A(n787), .ZN(n641) );
  NAND2_X1 U886 ( .A1(n763), .A2(n873), .ZN(n787) );
  INV_X1 U887 ( .A(n786), .ZN(n755) );
  NAND2_X1 U888 ( .A1(n760), .A2(n873), .ZN(n786) );
  INV_X1 U889 ( .A(n757), .ZN(n873) );
  AOI22_X1 U890 ( .A1(n3088gat), .A2(n3095gat), .B1(n3087gat), .B2(n3093gat), 
        .ZN(n757) );
  NOR2_X1 U891 ( .A1(n763), .A2(n872), .ZN(n760) );
  AOI21_X1 U892 ( .B1(n3087gat), .B2(n3095gat), .A(n667), .ZN(n872) );
  INV_X1 U893 ( .A(n583), .ZN(n667) );
  NAND2_X1 U894 ( .A1(n3093gat), .A2(n3086gat), .ZN(n583) );
  AOI21_X1 U895 ( .B1(n3086gat), .B2(n3095gat), .A(n668), .ZN(n763) );
  AND2_X1 U896 ( .A1(n3093gat), .A2(n3085gat), .ZN(n668) );
  NAND2_X1 U897 ( .A1(n874), .A2(n931gat), .ZN(n2709gat) );
  NAND2_X1 U898 ( .A1(n875), .A2(n557), .ZN(n2708gat) );
  NAND3_X1 U899 ( .A1(n876), .A2(n744), .A3(n877), .ZN(n2704gat) );
  OR3_X1 U900 ( .A1(n710), .A2(n3085gat), .A3(n709), .ZN(n744) );
  NAND3_X1 U901 ( .A1(n3088gat), .A2(n726), .A3(n723), .ZN(n709) );
  AND3_X1 U902 ( .A1(n584), .A2(n510), .A3(n3093gat), .ZN(n723) );
  INV_X1 U903 ( .A(n3087gat), .ZN(n726) );
  INV_X1 U904 ( .A(n3086gat), .ZN(n710) );
  NAND3_X1 U905 ( .A1(n713), .A2(n580), .A3(n585), .ZN(n876) );
  INV_X1 U906 ( .A(n712), .ZN(n585) );
  NAND3_X1 U907 ( .A1(n3087gat), .A2(n510), .A3(n665), .ZN(n712) );
  INV_X1 U908 ( .A(n3088gat), .ZN(n580) );
  NAND3_X1 U909 ( .A1(n3086gat), .A2(n510), .A3(n665), .ZN(n713) );
  AND3_X1 U910 ( .A1(n584), .A2(n749), .A3(n3095gat), .ZN(n665) );
  INV_X1 U911 ( .A(n3085gat), .ZN(n749) );
  NOR2_X1 U912 ( .A1(n3083gat), .A2(n3084gat), .ZN(n584) );
  NAND2_X1 U913 ( .A1(n530), .A2(n878), .ZN(n2702gat) );
  NAND2_X1 U914 ( .A1(n879), .A2(n531), .ZN(n2693gat) );
  OAI21_X1 U915 ( .B1(n2454gat), .B2(n544), .A(n880), .ZN(n2684gat) );
  XNOR2_X1 U916 ( .A(n881), .B(n882), .ZN(n2646gat) );
  XOR2_X1 U917 ( .A(n992), .B(n3128gat), .Z(n882) );
  XOR2_X1 U918 ( .A(n2339gat), .B(n3127gat), .Z(n881) );
  XNOR2_X1 U919 ( .A(n883), .B(n884), .ZN(n2613gat) );
  XNOR2_X1 U920 ( .A(n538), .B(n885), .ZN(n884) );
  XNOR2_X1 U921 ( .A(n993), .B(n527), .ZN(n885) );
  XNOR2_X1 U922 ( .A(n65), .B(n886), .ZN(n883) );
  XNOR2_X1 U923 ( .A(n67), .B(n512), .ZN(n886) );
  XNOR2_X1 U924 ( .A(n887), .B(n888), .ZN(n2579gat) );
  AOI21_X1 U925 ( .B1(n889), .B2(n64), .A(n890), .ZN(n888) );
  MUX2_X1 U926 ( .A(n891), .B(n823), .S(n53), .Z(n890) );
  NOR2_X1 U927 ( .A1(n62), .A2(n64), .ZN(n823) );
  NOR2_X1 U928 ( .A1(n64), .A2(n508), .ZN(n891) );
  XNOR2_X1 U929 ( .A(n62), .B(n53), .ZN(n889) );
  MUX2_X1 U930 ( .A(n892), .B(n893), .S(n84), .Z(n887) );
  NAND2_X1 U931 ( .A1(n742), .A2(n813), .ZN(n893) );
  NAND2_X1 U932 ( .A1(n57), .A2(n506), .ZN(n742) );
  OAI21_X1 U933 ( .B1(n524), .B2(n506), .A(n812), .ZN(n892) );
  NOR2_X1 U934 ( .A1(n746), .A2(n894), .ZN(n2556gat) );
  AOI21_X1 U935 ( .B1(n591), .B2(n509), .A(n498), .ZN(n746) );
  AND2_X1 U936 ( .A1(n747), .A2(n18), .ZN(n2436gat) );
  XNOR2_X1 U937 ( .A(n895), .B(n528), .ZN(n747) );
  NOR2_X1 U938 ( .A1(n896), .A2(n875), .ZN(n2396gat) );
  XNOR2_X1 U939 ( .A(n2403gat), .B(n897), .ZN(n875) );
  NOR2_X1 U940 ( .A1(n894), .A2(n880), .ZN(n2387gat) );
  NAND2_X1 U941 ( .A1(n898), .A2(n899), .ZN(n880) );
  OAI21_X1 U942 ( .B1(n1899gat), .B2(n2139gat), .A(n526), .ZN(n899) );
  INV_X1 U943 ( .A(n895), .ZN(n898) );
  NOR2_X1 U944 ( .A1(n877), .A2(n894), .ZN(n2330gat) );
  NOR2_X1 U945 ( .A1(n874), .A2(n896), .ZN(n2198gat) );
  NOR2_X1 U946 ( .A1(n752), .A2(n896), .ZN(n2197gat) );
  XNOR2_X1 U947 ( .A(n1003), .B(n594), .ZN(n752) );
  INV_X1 U948 ( .A(n900), .ZN(n594) );
  NOR2_X1 U949 ( .A1(n896), .A2(n751), .ZN(n2196gat) );
  OAI21_X1 U950 ( .B1(n901), .B2(n522), .A(n900), .ZN(n751) );
  NAND2_X1 U951 ( .A1(n901), .A2(n522), .ZN(n900) );
  NOR2_X1 U952 ( .A1(n897), .A2(n2403gat), .ZN(n901) );
  NOR2_X1 U953 ( .A1(n879), .A2(n902), .ZN(n2194gat) );
  AND2_X1 U954 ( .A1(n2262gat), .A2(n518), .ZN(n879) );
  AND4_X1 U955 ( .A1(n545), .A2(n903), .A3(n577), .A4(n1312gat), .ZN(n2163gat)
         );
  NOR2_X1 U956 ( .A1(n902), .A2(n878), .ZN(n2057gat) );
  NAND2_X1 U957 ( .A1(n904), .A2(n905), .ZN(n878) );
  OAI21_X1 U958 ( .B1(n2262gat), .B2(n518), .A(n550), .ZN(n905) );
  INV_X1 U959 ( .A(n628), .ZN(n904) );
  NOR3_X1 U960 ( .A1(n518), .A2(n2262gat), .A3(n550), .ZN(n628) );
  NOR2_X1 U961 ( .A1(n610), .A2(n906), .ZN(n2017gat) );
  NOR3_X1 U962 ( .A1(n2040gat), .A2(n1775gat), .A3(n1316gat), .ZN(n2015gat) );
  NOR2_X1 U963 ( .A1(n906), .A2(n907), .ZN(n1927gat) );
  NOR2_X1 U964 ( .A1(n908), .A2(n909), .ZN(n1915gat) );
  INV_X1 U965 ( .A(n498), .ZN(n908) );
  INV_X1 U966 ( .A(n896), .ZN(n19) );
  NAND2_X1 U967 ( .A1(n625), .A2(n20), .ZN(n896) );
  MUX2_X1 U968 ( .A(n910), .B(n911), .S(n2989gat), .Z(n625) );
  NAND2_X1 U969 ( .A1(n912), .A2(n913), .ZN(n910) );
  NOR3_X1 U970 ( .A1(n914), .A2(n1001), .A3(n1002), .ZN(n1882gat) );
  INV_X1 U971 ( .A(n915), .ZN(n914) );
  NOR2_X1 U972 ( .A1(n3099gat), .A2(n31), .ZN(n1827gat) );
  NOR2_X1 U973 ( .A1(n907), .A2(n909), .ZN(n1800gat) );
  NAND3_X1 U974 ( .A1(n514), .A2(n548), .A3(n913), .ZN(n909) );
  NOR3_X1 U975 ( .A1(n2347gat), .A2(n2440gat), .A3(n505), .ZN(n913) );
  INV_X1 U976 ( .A(n894), .ZN(n18) );
  NAND2_X1 U977 ( .A1(n626), .A2(n20), .ZN(n894) );
  INV_X1 U978 ( .A(n902), .ZN(n20) );
  OAI211_X1 U979 ( .C1(n998), .C2(n610), .A(n577), .B(n916), .ZN(n902) );
  AND2_X1 U980 ( .A1(n2037gat), .A2(n2095gat), .ZN(n916) );
  NAND2_X1 U981 ( .A1(n917), .A2(n496), .ZN(n577) );
  NAND4_X1 U982 ( .A1(n2506gat), .A2(n2502gat), .A3(n918), .A4(n2658gat), .ZN(
        n496) );
  NOR2_X1 U983 ( .A1(n999), .A2(n1000), .ZN(n918) );
  AND2_X1 U984 ( .A1(n2021gat), .A2(n533), .ZN(n610) );
  AND3_X1 U985 ( .A1(n919), .A2(n920), .A3(n921), .ZN(n626) );
  MUX2_X1 U986 ( .A(n922), .B(n923), .S(n994), .Z(n921) );
  NAND2_X1 U987 ( .A1(n498), .A2(n2989gat), .ZN(n922) );
  NOR2_X1 U988 ( .A1(n591), .A2(n509), .ZN(n498) );
  NAND2_X1 U989 ( .A1(n96), .A2(n895), .ZN(n591) );
  INV_X1 U990 ( .A(n924), .ZN(n920) );
  AOI211_X1 U991 ( .C1(n996), .C2(n995), .A(n2989gat), .B(n907), .ZN(n924) );
  NAND4_X1 U992 ( .A1(n500), .A2(n995), .A3(n996), .A4(n925), .ZN(n919) );
  NOR4_X1 U993 ( .A1(n526), .A2(n588), .A3(n513), .A4(n1899gat), .ZN(n500) );
  NOR2_X1 U994 ( .A1(n926), .A2(n927), .ZN(n1793gat) );
  INV_X1 U995 ( .A(n928), .ZN(n926) );
  NOR2_X1 U996 ( .A1(n3106gat), .A2(n602), .ZN(n1745gat) );
  AND2_X1 U997 ( .A1(n1775gat), .A2(n1771gat), .ZN(n602) );
  NOR4_X1 U998 ( .A1(n603), .A2(n508), .A3(n929), .A4(n930), .ZN(n1721gat) );
  INV_X1 U999 ( .A(n738), .ZN(n929) );
  NOR2_X1 U1000 ( .A1(n813), .A2(n53), .ZN(n738) );
  NAND2_X1 U1001 ( .A1(n63), .A2(n524), .ZN(n813) );
  NOR2_X1 U1002 ( .A1(n681), .A2(n675), .ZN(n603) );
  AND3_X1 U1003 ( .A1(n931), .A2(n504), .A3(n851), .ZN(n675) );
  AND4_X1 U1004 ( .A1(n741), .A2(n543), .A3(n507), .A4(n504), .ZN(n681) );
  NOR2_X1 U1005 ( .A1(n932), .A2(n599), .ZN(n1696gat) );
  NOR4_X1 U1006 ( .A1(n925), .A2(n509), .A3(n933), .A4(n528), .ZN(n1636gat) );
  INV_X1 U1007 ( .A(n2989gat), .ZN(n925) );
  NOR4_X1 U1008 ( .A1(n1006), .A2(n1007), .A3(n523), .A4(n507), .ZN(n1620gat)
         );
  NOR2_X1 U1009 ( .A1(n932), .A2(n597), .ZN(n1613gat) );
  NOR2_X1 U1010 ( .A1(n932), .A2(n934), .ZN(n1610gat) );
  INV_X1 U1011 ( .A(n1606gat), .ZN(n934) );
  OAI211_X1 U1012 ( .C1(n32), .C2(n546), .A(n915), .B(n2472gat), .ZN(n932) );
  NAND2_X1 U1013 ( .A1(n917), .A2(n2830gat), .ZN(n915) );
  NAND2_X1 U1014 ( .A1(n2446gat), .A2(n2450gat), .ZN(n2830gat) );
  INV_X1 U1015 ( .A(n3100gat), .ZN(n917) );
  NOR2_X1 U1016 ( .A1(n2454gat), .A2(n271gat), .ZN(n1606gat) );
  AND3_X1 U1017 ( .A1(n1312gat), .A2(n935), .A3(n936), .ZN(n1593gat) );
  NOR2_X1 U1018 ( .A1(n927), .A2(n575), .ZN(n1567gat) );
  NAND3_X1 U1019 ( .A1(n935), .A2(n877), .A3(n97), .ZN(n575) );
  NOR2_X1 U1020 ( .A1(n513), .A2(n532), .ZN(n877) );
  NOR4_X1 U1021 ( .A1(n1899gat), .A2(n588), .A3(n587), .A4(n927), .ZN(n1565gat) );
  NAND3_X1 U1022 ( .A1(n2440gat), .A2(n522), .A3(n937), .ZN(n927) );
  NOR3_X1 U1023 ( .A1(n2394gat), .A2(n1003), .A3(n2403gat), .ZN(n937) );
  NAND2_X1 U1024 ( .A1(n513), .A2(n526), .ZN(n587) );
  NOR3_X1 U1025 ( .A1(n923), .A2(n906), .A3(n938), .ZN(n1564gat) );
  INV_X1 U1026 ( .A(n911), .ZN(n938) );
  NAND4_X1 U1027 ( .A1(n912), .A2(n2440gat), .A3(n522), .A4(n505), .ZN(n911)
         );
  INV_X1 U1028 ( .A(n903), .ZN(n906) );
  NAND4_X1 U1029 ( .A1(n939), .A2(n1003), .A3(n928), .A4(n3149gat), .ZN(n903)
         );
  NAND3_X1 U1030 ( .A1(n1767gat), .A2(n1834gat), .A3(n533), .ZN(n3149gat) );
  OAI21_X1 U1031 ( .B1(n2989gat), .B2(n907), .A(n923), .ZN(n928) );
  NAND2_X1 U1032 ( .A1(n895), .A2(n935), .ZN(n907) );
  NOR3_X1 U1033 ( .A1(n1899gat), .A2(n2139gat), .A3(n526), .ZN(n895) );
  MUX2_X1 U1034 ( .A(n940), .B(n941), .S(n514), .Z(n939) );
  NOR3_X1 U1035 ( .A1(n942), .A2(n522), .A3(n858), .ZN(n941) );
  INV_X1 U1036 ( .A(n931), .ZN(n858) );
  MUX2_X1 U1037 ( .A(n943), .B(n944), .S(n945), .Z(n942) );
  OR2_X1 U1038 ( .A1(n505), .A2(n946), .ZN(n944) );
  MUX2_X1 U1039 ( .A(n947), .B(n897), .S(n741), .Z(n943) );
  NAND2_X1 U1040 ( .A1(n505), .A2(n529), .ZN(n897) );
  NAND2_X1 U1041 ( .A1(n2440gat), .A2(n505), .ZN(n947) );
  MUX2_X1 U1042 ( .A(n948), .B(n874), .S(n522), .Z(n940) );
  NOR3_X1 U1043 ( .A1(n949), .A2(n931), .A3(n946), .ZN(n948) );
  XOR2_X1 U1044 ( .A(n741), .B(n529), .Z(n946) );
  NOR2_X1 U1045 ( .A1(n511), .A2(n523), .ZN(n741) );
  NOR2_X1 U1046 ( .A1(n523), .A2(n402gat), .ZN(n931) );
  MUX2_X1 U1047 ( .A(n950), .B(n945), .S(n505), .Z(n949) );
  NAND2_X1 U1048 ( .A1(n398gat), .A2(n945), .ZN(n950) );
  NAND4_X1 U1049 ( .A1(n936), .A2(n2989gat), .A3(n509), .A4(n528), .ZN(n923)
         );
  OAI21_X1 U1050 ( .B1(n533), .B2(n1763gat), .A(n2102gat), .ZN(n2989gat) );
  NOR4_X1 U1051 ( .A1(n951), .A2(n522), .A3(n588), .A4(n933), .ZN(n1516gat) );
  INV_X1 U1052 ( .A(n936), .ZN(n933) );
  NOR3_X1 U1053 ( .A1(n1899gat), .A2(n97), .A3(n513), .ZN(n936) );
  INV_X1 U1054 ( .A(n935), .ZN(n588) );
  NOR2_X1 U1055 ( .A1(n509), .A2(n96), .ZN(n935) );
  NAND2_X1 U1056 ( .A1(n874), .A2(n912), .ZN(n951) );
  NOR2_X1 U1057 ( .A1(n548), .A2(n514), .ZN(n912) );
  NOR2_X1 U1058 ( .A1(n505), .A2(n529), .ZN(n874) );
  INV_X1 U1059 ( .A(n599), .ZN(n15) );
  NAND3_X1 U1060 ( .A1(n852), .A2(n507), .A3(n851), .ZN(n599) );
  NOR2_X1 U1061 ( .A1(n1007), .A2(n2454gat), .ZN(n851) );
  NOR3_X1 U1062 ( .A1(n930), .A2(n62), .A3(n952), .ZN(n1391gat) );
  INV_X1 U1063 ( .A(n809), .ZN(n952) );
  NOR2_X1 U1064 ( .A1(n812), .A2(n53), .ZN(n809) );
  NAND2_X1 U1065 ( .A1(n524), .A2(n506), .ZN(n812) );
  NAND4_X1 U1066 ( .A1(n64), .A2(n512), .A3(n65), .A4(n953), .ZN(n930) );
  NOR3_X1 U1067 ( .A1(n67), .A2(n69), .A3(n68), .ZN(n953) );
  INV_X1 U1068 ( .A(n597), .ZN(n13) );
  NAND2_X1 U1069 ( .A1(n853), .A2(n507), .ZN(n597) );
  NOR3_X1 U1070 ( .A1(n511), .A2(n2454gat), .A3(n945), .ZN(n853) );
  INV_X1 U1071 ( .A(n852), .ZN(n945) );
  NOR2_X1 U1072 ( .A1(n504), .A2(n523), .ZN(n852) );
  XNOR2_X1 U1073 ( .A(n954), .B(n955), .ZN(n1269gat) );
  XOR2_X1 U1074 ( .A(n956), .B(n957), .Z(n955) );
  XNOR2_X1 U1075 ( .A(n531), .B(n1005), .ZN(n957) );
  XNOR2_X1 U1076 ( .A(n530), .B(n1004), .ZN(n956) );
  XOR2_X1 U1077 ( .A(n958), .B(n959), .Z(n954) );
  XNOR2_X1 U1078 ( .A(n539), .B(n931gat), .ZN(n959) );
  XNOR2_X1 U1079 ( .A(n75), .B(n76), .ZN(n958) );
  INV_X1 U1080 ( .A(blif_reset_net), .ZN(n1) );
  SDFFS_X2 n673gat_reg ( .D(n2897gat), .SI(n667gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n562), .Q(n673gat), .QN(n525) );
  SDFFS_X2 n398gat_reg ( .D(n3069gat), .SI(n17), .SE(test_se), .CK(
        blif_clk_net), .SN(n563), .Q(n398gat), .QN(n523) );
  SDFFS_X2 n402gat_reg ( .D(n3070gat), .SI(n398gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n561), .Q(n402gat), .QN(n507) );
  SDFFS_X2 n919gat_reg ( .D(n3072gat), .SI(n21), .SE(test_se), .CK(
        blif_clk_net), .SN(n561), .Q(n511), .QN(n1007) );
  SDFFS_X2 n846gat_reg ( .D(n3071gat), .SI(n119), .SE(test_se), .CK(
        blif_clk_net), .SN(n562), .Q(n504), .QN(n1006) );
  SDFFS_X2 n2510gat_reg ( .D(n748gat), .SI(n2506gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n561), .Q(n121), .QN(n999) );
  SDFFS_X2 n271gat_reg ( .D(n3065gat), .SI(n10), .SE(test_se), .CK(
        blif_clk_net), .SN(n562), .Q(n271gat), .QN(n517) );
  SDFFS_X2 n160gat_reg ( .D(n3067gat), .SI(n12), .SE(test_se), .CK(
        blif_clk_net), .SN(n562), .Q(n120), .QN(n25) );
  SDFFS_X2 n337gat_reg ( .D(n3066gat), .SI(n977), .SE(test_se), .CK(
        blif_clk_net), .SN(n561), .Q(n544), .QN(n991) );
  SDFFS_X2 n842gat_reg ( .D(n3073gat), .SI(n838gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n559), .Q(n119), .QN(n516) );
  SDFFS_X2 n341gat_reg ( .D(n3068gat), .SI(n544), .SE(test_se), .CK(
        blif_clk_net), .SN(n561), .Q(n341gat), .QN(n519) );
  SDFFS_X2 n2522gat_reg ( .D(n55gat), .SI(n44), .SE(test_se), .CK(blif_clk_net), .SN(n561), .Q(n118), .QN(n965) );
  SDFFS_X2 n2472gat_reg ( .D(n1620gat), .SI(n102), .SE(test_se), .CK(
        blif_clk_net), .SN(n561), .Q(n2472gat), .QN(n30) );
  SDFFS_X2 n2319gat_reg ( .D(n30), .SI(n93), .SE(test_se), .CK(blif_clk_net), 
        .SN(n559), .Q(n117), .QN(n31) );
  SDFFS_X2 n1821gat_reg ( .D(n1827gat), .SI(n1807gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n559), .Q(n115), .QN(n32) );
  SDFFS_X2 n2029gat_reg ( .D(n32), .SI(n23), .SE(test_se), .CK(blif_clk_net), 
        .SN(n560), .Q(n111), .QN(n33) );
  SDFFS_X2 n1829gat_reg ( .D(n33), .SI(n115), .SE(test_se), .CK(blif_clk_net), 
        .SN(n562), .Q(n546) );
  SDFFS_X2 n2476gat_reg ( .D(n55gat), .SI(n2472gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n561), .Q(n108), .QN(n970) );
  SDFFS_X2 n1068gat_reg ( .D(n2914gat), .SI(n539), .SE(test_se), .CK(
        blif_clk_net), .SN(n561), .Q(n107), .QN(n34) );
  SDFFS_X2 n957gat_reg ( .D(n2928gat), .SI(n931gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n562), .Q(n106), .QN(n515) );
  SDFFS_X2 n861gat_reg ( .D(n2927gat), .SI(n504), .SE(test_se), .CK(
        blif_clk_net), .SN(n561), .Q(n537), .QN(n990) );
  SDFFS_X2 n1294gat_reg ( .D(n2896gat), .SI(n531), .SE(test_se), .CK(
        blif_clk_net), .SN(n561), .Q(n105), .QN(n985) );
  SDFFS_X2 n1241gat_reg ( .D(n2922gat), .SI(n556), .SE(test_se), .CK(
        blif_clk_net), .SN(n560), .Q(n104), .QN(n980) );
  SDFFS_X2 n865gat_reg ( .D(n2894gat), .SI(n537), .SE(test_se), .CK(
        blif_clk_net), .SN(n560), .Q(n865gat) );
  SDFFS_X2 n1080gat_reg ( .D(n2921gat), .SI(n554), .SE(test_se), .CK(
        blif_clk_net), .SN(n562), .Q(n103), .QN(n37) );
  SDFFS_X2 n1148gat_reg ( .D(n2895gat), .SI(n530), .SE(test_se), .CK(
        blif_clk_net), .SN(n561), .Q(n535), .QN(n983) );
  SDFFS_X2 n2468gat_reg ( .D(n933gat), .SI(n14), .SE(test_se), .CK(
        blif_clk_net), .SN(n562), .Q(n102), .QN(n969) );
  SDFFS_X2 n2450gat_reg ( .D(1'b0), .SI(n2446gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n566), .Q(n2450gat), .QN(n3148gat) );
  SDFFS_X2 n148gat_reg ( .D(n38), .SI(test_si1), .SE(test_se), .CK(
        blif_clk_net), .SN(n566), .Q(n148gat) );
  SDFFS_X2 n834gat_reg ( .D(n2923gat), .SI(n830gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n566), .Q(n834gat), .QN(n38) );
  SDFFS_X2 n2526gat_reg ( .D(n504gat), .SI(n118), .SE(test_se), .CK(
        blif_clk_net), .SN(n566), .Q(n101), .QN(n966) );
  SDFFS_X2 n2588gat_reg ( .D(n3016gat), .SI(n506), .SE(test_se), .CK(
        blif_clk_net), .SN(n563), .Q(n100), .QN(n1000) );
  SDFFS_X2 n2446gat_reg ( .D(n496), .SI(n2440gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n562), .Q(n2446gat) );
  SDFFS_X2 n1871gat_reg ( .D(n7), .SI(n55), .SE(test_se), .CK(blif_clk_net), 
        .SN(n565), .Q(n510), .QN(n3106gat) );
  SDFFS_X2 n2095gat_reg ( .D(n502), .SI(n60), .SE(test_se), .CK(blif_clk_net), 
        .SN(n566), .Q(n2095gat), .QN(n128) );
  SDFFS_X2 n2176gat_reg ( .D(n128), .SI(n98), .SE(test_se), .CK(blif_clk_net), 
        .SN(n566), .Q(n99), .QN(n129) );
  SDFFS_X2 n2169gat_reg ( .D(n129), .SI(n77), .SE(test_se), .CK(blif_clk_net), 
        .SN(n567), .Q(n98), .QN(n545) );
  SDFFS_X2 n2390gat_reg ( .D(n20), .SI(n2347gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n562), .Q(n95), .QN(n3128gat) );
  SDFFS_X2 n2262gat_reg ( .D(n3128gat), .SI(n534), .SE(test_se), .CK(
        blif_clk_net), .SN(n563), .Q(n2262gat) );
  SDFFS_X2 n2270gat_reg ( .D(n2194gat), .SI(n92), .SE(test_se), .CK(
        blif_clk_net), .SN(n562), .Q(n93), .QN(n3127gat) );
  SDFFS_X2 n2190gat_reg ( .D(n3127gat), .SI(n24), .SE(test_se), .CK(
        blif_clk_net), .SN(n563), .Q(n518), .QN(n997) );
  SDFFS_X2 n2495gat_reg ( .D(n493), .SI(n512), .SE(test_se), .CK(blif_clk_net), 
        .SN(n559), .Q(n992), .QN(n85) );
  SDFFS_X2 n2266gat_reg ( .D(n85), .SI(n2262gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n563), .Q(n92), .QN(n961) );
  SDFFS_X2 n2339gat_reg ( .D(n2057gat), .SI(n117), .SE(test_se), .CK(
        blif_clk_net), .SN(n563), .Q(n2339gat), .QN(n3126gat) );
  SDFFS_X2 n2135gat_reg ( .D(n3126gat), .SI(n1002), .SE(test_se), .CK(
        blif_clk_net), .SN(n563), .Q(n550) );
  SDFFS_X2 n1433gat_reg ( .D(n2983gat), .SI(n1394gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n560), .Q(n91), .QN(n112) );
  SDFFS_X2 n1316gat_reg ( .D(n112), .SI(n1312gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n563), .Q(n1316gat), .QN(n113) );
  SDFFS_X2 n1363gat_reg ( .D(n113), .SI(n521), .SE(test_se), .CK(blif_clk_net), 
        .SN(n559), .Q(n90), .QN(n114) );
  SDFFS_X2 n1312gat_reg ( .D(n114), .SI(n105), .SE(test_se), .CK(blif_clk_net), 
        .SN(n563), .Q(n1312gat) );
  SDFFS_X2 n2044gat_reg ( .D(n2015gat), .SI(n2040gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n559), .Q(n88), .QN(n132) );
  SDFFS_X2 n2037gat_reg ( .D(n132), .SI(n2033gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n572), .Q(n2037gat), .QN(n133) );
  SDFFS_X2 n2033gat_reg ( .D(n133), .SI(n111), .SE(test_se), .CK(blif_clk_net), 
        .SN(n572), .Q(n2033gat), .QN(n135) );
  SDFFS_X2 n2110gat_reg ( .D(n135), .SI(n2102gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n559), .Q(n87), .QN(n136) );
  SDFFS_X2 n2125gat_reg ( .D(n136), .SI(n86), .SE(test_se), .CK(blif_clk_net), 
        .SN(n559), .Q(n1002), .QN(n137) );
  SDFFS_X2 n2121gat_reg ( .D(n137), .SI(n78), .SE(test_se), .CK(blif_clk_net), 
        .SN(n559), .Q(n86), .QN(n138) );
  SDFFS_X2 n2117gat_reg ( .D(n138), .SI(n87), .SE(test_se), .CK(blif_clk_net), 
        .SN(n572), .Q(n78), .QN(n1001) );
  SDFFS_X2 n1880gat_reg ( .D(n1882gat), .SI(n510), .SE(test_se), .CK(
        blif_clk_net), .SN(n563), .Q(n533) );
  SDFFS_X2 n2155gat_reg ( .D(n2989gat), .SI(n528), .SE(test_se), .CK(
        blif_clk_net), .SN(n565), .Q(n77), .QN(n74) );
  SDFFS_X2 n2562gat_reg ( .D(n19), .SI(n527), .SE(test_se), .CK(blif_clk_net), 
        .SN(n564), .Q(n506), .QN(n63) );
  SDFFS_X2 n2440gat_reg ( .D(n63), .SI(n548), .SE(test_se), .CK(blif_clk_net), 
        .SN(n564), .Q(n2440gat), .QN(n529) );
  SDFFS_X2 n2343gat_reg ( .D(n2198gat), .SI(n2339gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n564), .Q(n524), .QN(n57) );
  SDFFS_X2 n2394gat_reg ( .D(n57), .SI(n95), .SE(test_se), .CK(blif_clk_net), 
        .SN(n564), .Q(n2394gat), .QN(n505) );
  SDFFS_X2 n2399gat_reg ( .D(n2396gat), .SI(n2394gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n564), .Q(n73), .QN(n53) );
  SDFFS_X2 n2403gat_reg ( .D(n53), .SI(n73), .SE(test_se), .CK(blif_clk_net), 
        .SN(n564), .Q(n2403gat), .QN(n514) );
  SDFFS_X2 n2203gat_reg ( .D(n2196gat), .SI(n518), .SE(test_se), .CK(
        blif_clk_net), .SN(n564), .Q(n508), .QN(n62) );
  SDFFS_X2 n2347gat_reg ( .D(n62), .SI(n524), .SE(test_se), .CK(blif_clk_net), 
        .SN(n564), .Q(n2347gat), .QN(n522) );
  SDFFS_X2 n2640gat_reg ( .D(n494), .SI(n993), .SE(test_se), .CK(blif_clk_net), 
        .SN(n564), .Q(n72), .QN(n84) );
  SDFFS_X2 n2644gat_reg ( .D(n84), .SI(n72), .SE(test_se), .CK(blif_clk_net), 
        .SN(n565), .Q(n71), .QN(n962) );
  SDFFS_X2 n2207gat_reg ( .D(n2197gat), .SI(n508), .SE(test_se), .CK(
        blif_clk_net), .SN(n565), .Q(n534), .QN(n64) );
  SDFFS_X2 n2407gat_reg ( .D(n64), .SI(n2403gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n564), .Q(n548), .QN(n1003) );
  SDFFS_X2 n2658gat_reg ( .D(n2579gat), .SI(n71), .SE(test_se), .CK(
        blif_clk_net), .SN(n565), .Q(n2658gat) );
  SDFFS_X2 n1389gat_reg ( .D(n1793gat), .SI(n90), .SE(test_se), .CK(
        blif_clk_net), .SN(n571), .Q(n70), .QN(n981) );
  SDFFS_X2 n2454gat_reg ( .D(n2163gat), .SI(n2450gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n564), .Q(n2454gat), .QN(n543) );
  SDFFS_X2 n1767gat_reg ( .D(n15), .SI(n1763gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n565), .Q(n1767gat) );
  SDFFS_X2 n1775gat_reg ( .D(n1696gat), .SI(n1771gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n565), .Q(n1775gat), .QN(n116) );
  SDFFS_X2 n2592gat_reg ( .D(n116), .SI(n100), .SE(test_se), .CK(blif_clk_net), 
        .SN(n560), .Q(n2592gat), .QN(n123) );
  SDFFS_X2 n2179gat_reg ( .D(n492), .SI(n99), .SE(test_se), .CK(blif_clk_net), 
        .SN(n567), .Q(n61), .QN(n972) );
  SDFFS_X2 n2091gat_reg ( .D(n491), .SI(n26), .SE(test_se), .CK(blif_clk_net), 
        .SN(n568), .Q(n60), .QN(n996) );
  SDFFS_X2 n2626gat_reg ( .D(n18), .SI(n58), .SE(test_se), .CK(blif_clk_net), 
        .SN(n568), .Q(n59), .QN(n65) );
  SDFFS_X2 n1899gat_reg ( .D(n65), .SI(n533), .SE(test_se), .CK(blif_clk_net), 
        .SN(n568), .Q(n1899gat), .QN(n532) );
  SDFFS_X2 n2490gat_reg ( .D(n2330gat), .SI(n108), .SE(test_se), .CK(
        blif_clk_net), .SN(n568), .Q(n512), .QN(n66) );
  SDFFS_X2 n2139gat_reg ( .D(n66), .SI(n550), .SE(test_se), .CK(blif_clk_net), 
        .SN(n568), .Q(n2139gat), .QN(n513) );
  SDFFS_X2 n2622gat_reg ( .D(n2387gat), .SI(n27), .SE(test_se), .CK(
        blif_clk_net), .SN(n568), .Q(n58), .QN(n67) );
  SDFFS_X2 n2061gat_reg ( .D(n67), .SI(n88), .SE(test_se), .CK(blif_clk_net), 
        .SN(n568), .Q(n526), .QN(n97) );
  SDFFS_X2 n2543gat_reg ( .D(n2436gat), .SI(n101), .SE(test_se), .CK(
        blif_clk_net), .SN(n568), .Q(n527), .QN(n69) );
  SDFFS_X2 n2143gat_reg ( .D(n69), .SI(n2139gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n568), .Q(n528), .QN(n96) );
  SDFFS_X2 n2634gat_reg ( .D(n495), .SI(n538), .SE(test_se), .CK(blif_clk_net), 
        .SN(n560), .Q(n993), .QN(n89) );
  SDFFS_X2 n1975gat_reg ( .D(n89), .SI(n1899gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n568), .Q(n56), .QN(n963) );
  SDFFS_X2 n2630gat_reg ( .D(n2556gat), .SI(n59), .SE(test_se), .CK(
        blif_clk_net), .SN(n568), .Q(n538), .QN(n68) );
  SDFFS_X2 n1850gat_reg ( .D(n68), .SI(n1834gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n570), .Q(n55), .QN(n509) );
  SDFFS_X2 n1332gat_reg ( .D(n1565gat), .SI(n1316gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n559), .Q(n54), .QN(n110) );
  SDFFS_X2 n1740gat_reg ( .D(n110), .SI(n1678gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n570), .Q(n52), .QN(n994) );
  SDFFS_X2 n1678gat_reg ( .D(n94), .SI(n8), .SE(test_se), .CK(blif_clk_net), 
        .SN(n571), .Q(n1678gat) );
  SDFFS_X2 n1508gat_reg ( .D(n1636gat), .SI(n51), .SE(test_se), .CK(
        blif_clk_net), .SN(n559), .Q(n982) );
  SDFFS_X2 n1394gat_reg ( .D(n1516gat), .SI(n70), .SE(test_se), .CK(
        blif_clk_net), .SN(n560), .Q(n1394gat), .QN(n109) );
  SDFFS_X2 n1496gat_reg ( .D(n109), .SI(n555), .SE(test_se), .CK(blif_clk_net), 
        .SN(n570), .Q(n51), .QN(n995) );
  SDFFS_X2 n2506gat_reg ( .D(n2613gat), .SI(n2502gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n568), .Q(n2506gat) );
  SDFFS_X2 n1121gat_reg ( .D(n2952gat), .SI(n103), .SE(test_se), .CK(
        blif_clk_net), .SN(n570), .Q(n557), .QN(n76) );
  SDFFS_X2 n1072gat_reg ( .D(n2919gat), .SI(n107), .SE(test_se), .CK(
        blif_clk_net), .SN(n570), .Q(n554), .QN(n1005) );
  SDFFS_X2 n1035gat_reg ( .D(n2918gat), .SI(n106), .SE(test_se), .CK(
        blif_clk_net), .SN(n570), .Q(n558), .QN(n75) );
  SDFFS_X2 n777gat_reg ( .D(n2915gat), .SI(n11), .SE(test_se), .CK(
        blif_clk_net), .SN(n570), .Q(n45), .QN(n80) );
  SDFFS_X2 n1135gat_reg ( .D(n2912gat), .SI(n557), .SE(test_se), .CK(
        blif_clk_net), .SN(n570), .Q(n530) );
  SDFFS_X2 n931gat_reg ( .D(n2911gat), .SI(n511), .SE(test_se), .CK(
        blif_clk_net), .SN(n570), .Q(n931gat), .QN(n551) );
  SDFFS_X2 n1282gat_reg ( .D(n2910gat), .SI(n104), .SE(test_se), .CK(
        blif_clk_net), .SN(n569), .Q(n531) );
  SDFFS_X2 n1045gat_reg ( .D(n2909gat), .SI(n558), .SE(test_se), .CK(
        blif_clk_net), .SN(n569), .Q(n539) );
  SDFFS_X2 n1197gat_reg ( .D(n2908gat), .SI(n535), .SE(test_se), .CK(
        blif_clk_net), .SN(n569), .Q(n1197gat) );
  SDFFS_X2 n1226gat_reg ( .D(n2907gat), .SI(n1197gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n569), .Q(n556), .QN(n1004) );
  SDFFS_X2 n2518gat_reg ( .D(n2971gat), .SI(n549), .SE(test_se), .CK(
        blif_clk_net), .SN(n570), .Q(n44), .QN(n964) );
  SDFFS_X2 n667gat_reg ( .D(n2904gat), .SI(n35), .SE(test_se), .CK(
        blif_clk_net), .SN(n569), .Q(n667gat) );
  SDFFS_X2 n553gat_reg ( .D(n2903gat), .SI(n470gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n569), .Q(n43), .QN(n988) );
  SDFFS_X2 n561gat_reg ( .D(n2901gat), .SI(n43), .SE(test_se), .CK(
        blif_clk_net), .SN(n569), .Q(n36), .QN(n81) );
  SDFFS_X2 n659gat_reg ( .D(n2891gat), .SI(n614gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n569), .Q(n35), .QN(n79) );
  SDFFS_X2 n366gat_reg ( .D(n2890gat), .SI(n341gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n569), .Q(n29), .QN(n989) );
  SDFFS_X2 n322gat_reg ( .D(n2888gat), .SI(n541), .SE(test_se), .CK(
        blif_clk_net), .SN(n569), .Q(n28), .QN(n987) );
  SDFFS_X2 n318gat_reg ( .D(n2887gat), .SI(n520), .SE(test_se), .CK(
        blif_clk_net), .SN(n569), .Q(n541), .QN(n82) );
  SDFFS_X2 n314gat_reg ( .D(n2886gat), .SI(n271gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n569), .Q(n520), .QN(n83) );
  SDFFS_X2 n2599gat_reg ( .D(n3010gat), .SI(n2592gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n570), .Q(n27), .QN(n967) );
  SDFFS_X2 n2102gat_reg ( .D(n1606gat), .SI(n22), .SE(test_se), .CK(
        blif_clk_net), .SN(n564), .Q(n2102gat) );
  SDFFS_X2 n1763gat_reg ( .D(n1610gat), .SI(n1748gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n563), .Q(n1763gat) );
  SDFFS_X2 n1834gat_reg ( .D(n13), .SI(n546), .SE(test_se), .CK(blif_clk_net), 
        .SN(n571), .Q(n1834gat) );
  SDFFS_X2 n2084gat_reg ( .D(n3149gat), .SI(n526), .SE(test_se), .CK(
        blif_clk_net), .SN(n571), .Q(n26), .QN(n986) );
  SDFFS_X2 n2182gat_reg ( .D(n489), .SI(n61), .SE(test_se), .CK(blif_clk_net), 
        .SN(n572), .Q(n24), .QN(n971) );
  SDFFS_X2 n2040gat_reg ( .D(n6), .SI(n2037gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n572), .Q(n2040gat) );
  SDFFS_X2 n2021gat_reg ( .D(n488), .SI(n56), .SE(test_se), .CK(blif_clk_net), 
        .SN(n572), .Q(n2021gat) );
  SDFFS_X2 n2025gat_reg ( .D(n2017gat), .SI(n2021gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n559), .Q(n23), .QN(n134) );
  SDFFS_X2 n2099gat_reg ( .D(n134), .SI(n2095gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n562), .Q(n22), .QN(n998) );
  SDFFS_X2 n2502gat_reg ( .D(n2646gat), .SI(n992), .SE(test_se), .CK(
        blif_clk_net), .SN(n563), .Q(n2502gat) );
  SDFFS_X2 n816gat_reg ( .D(n2920gat), .SI(n45), .SE(test_se), .CK(
        blif_clk_net), .SN(n566), .Q(n816gat), .QN(n547) );
  SDFFS_X2 n680gat_reg ( .D(n2913gat), .SI(n673gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n566), .Q(n680gat), .QN(n540) );
  SDFFS_X2 n580gat_reg ( .D(n2905gat), .SI(n36), .SE(test_se), .CK(
        blif_clk_net), .SN(n566), .Q(n580gat), .QN(n552) );
  SDFFS_X2 n883gat_reg ( .D(n2929gat), .SI(n865gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n567), .Q(n21), .QN(n48) );
  SDFFS_X2 n388gat_reg ( .D(n48), .SI(n384gat), .SE(test_se), .CK(blif_clk_net), .SN(n567), .Q(n17), .QN(n978) );
  SDFFS_X2 n824gat_reg ( .D(n2900gat), .SI(n820gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n567), .Q(n824gat), .QN(n46) );
  SDFFS_X2 n331gat_reg ( .D(n46), .SI(n536), .SE(test_se), .CK(blif_clk_net), 
        .SN(n560), .Q(n977), .QN(n542) );
  SDFFS_X2 n684gat_reg ( .D(n2916gat), .SI(n680gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n560), .Q(n16), .QN(n49) );
  SDFFS_X2 n327gat_reg ( .D(n49), .SI(n28), .SE(test_se), .CK(blif_clk_net), 
        .SN(n567), .Q(n536), .QN(n976) );
  SDFFS_X2 n820gat_reg ( .D(n2925gat), .SI(n816gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n567), .Q(n820gat), .QN(n47) );
  SDFFS_X2 n463gat_reg ( .D(n47), .SI(n402gat), .SE(test_se), .CK(blif_clk_net), .SN(n567), .Q(n463gat) );
  SDFFS_X2 n699gat_reg ( .D(n2899gat), .SI(n16), .SE(test_se), .CK(
        blif_clk_net), .SN(n567), .Q(n699gat), .QN(n50) );
  SDFFS_X2 n384gat_reg ( .D(n50), .SI(n29), .SE(test_se), .CK(blif_clk_net), 
        .SN(n567), .Q(n384gat) );
  SDFFS_X2 n584gat_reg ( .D(n2898gat), .SI(n580gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n566), .Q(n553), .QN(n984) );
  SDFFS_X2 n2464gat_reg ( .D(n567gat), .SI(n9), .SE(test_se), .CK(blif_clk_net), .SN(n567), .Q(n14), .QN(n968) );
  SDFFS_X2 n614gat_reg ( .D(n2892gat), .SI(n553), .SE(test_se), .CK(
        blif_clk_net), .SN(n565), .Q(n614gat), .QN(n42) );
  SDFFS_X2 n156gat_reg ( .D(n42), .SI(n975), .SE(test_se), .CK(blif_clk_net), 
        .SN(n565), .Q(n12), .QN(n979) );
  SDFFS_X2 n707gat_reg ( .D(n2917gat), .SI(n699gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n565), .Q(n11), .QN(n39) );
  SDFFS_X2 n152gat_reg ( .D(n39), .SI(n148gat), .SE(test_se), .CK(blif_clk_net), .SN(n560), .Q(n975) );
  SDFFS_X2 n838gat_reg ( .D(n2924gat), .SI(n834gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n565), .Q(n838gat), .QN(n40) );
  SDFFS_X2 n256gat_reg ( .D(n40), .SI(n120), .SE(test_se), .CK(blif_clk_net), 
        .SN(n565), .Q(n10), .QN(n974) );
  SDFFS_X2 n830gat_reg ( .D(n2926gat), .SI(n824gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n566), .Q(n830gat), .QN(n41) );
  SDFFS_X2 n470gat_reg ( .D(n41), .SI(n463gat), .SE(test_se), .CK(blif_clk_net), .SN(n566), .Q(n470gat) );
  SDFFS_X2 n2458gat_reg ( .D(n123), .SI(n2454gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n560), .Q(n9), .QN(n141) );
  SDFFS_X2 n2514gat_reg ( .D(n141), .SI(n121), .SE(test_se), .CK(blif_clk_net), 
        .SN(n567), .Q(n549) );
  SDFFS_X2 n1771gat_reg ( .D(n1613gat), .SI(test_si2), .SE(test_se), .CK(
        blif_clk_net), .SN(n572), .Q(n1771gat) );
  SDFFS_X2 n1336gat_reg ( .D(n1391gat), .SI(n54), .SE(test_se), .CK(
        blif_clk_net), .SN(n570), .Q(n1336gat) );
  SDFFS_X2 n1748gat_reg ( .D(n1927gat), .SI(n52), .SE(test_se), .CK(
        blif_clk_net), .SN(n571), .Q(n1748gat) );
  SDFFS_X2 n1675gat_reg ( .D(n500), .SI(n1596gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n571), .Q(n8), .QN(n973) );
  SDFFS_X2 n1807gat_reg ( .D(n498), .SI(n1775gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n571), .Q(n1807gat) );
  SDFFS_X2 n1340gat_reg ( .D(n1567gat), .SI(n1336gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n571), .Q(n521), .QN(n142) );
  SDFFS_X2 n1456gat_reg ( .D(n1564gat), .SI(n91), .SE(test_se), .CK(
        blif_clk_net), .SN(n571), .Q(n1456gat) );
  SDFFS_X2 n1525gat_reg ( .D(n499), .SI(n982), .SE(test_se), .CK(blif_clk_net), 
        .SN(n571), .Q(n1525gat) );
  SDFFS_X2 n1462gat_reg ( .D(n1915gat), .SI(n1456gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n571), .Q(n555), .QN(n1008) );
  SDFFS_X2 n1596gat_reg ( .D(n1800gat), .SI(n5), .SE(test_se), .CK(
        blif_clk_net), .SN(n571), .Q(n1596gat) );
  SDFFS_X2 n1588gat_reg ( .D(n1593gat), .SI(n1525gat), .SE(test_se), .CK(
        blif_clk_net), .SN(n560), .Q(n5), .QN(n960) );
endmodule

