
module multdiv ( data_operandA, data_operandB, ctrl_MULT, ctrl_DIV, clock, 
        data_result, data_exception, data_resultRDY );
  input [31:0] data_operandA;
  input [31:0] data_operandB;
  output [31:0] data_result;
  input ctrl_MULT, ctrl_DIV, clock;
  output data_exception, data_resultRDY;
  wire   nop, shift, op_mult, op_div, div_ready, n_1_net__31_, n_1_net__22_,
         n_1_net__21_, n_1_net__20_, n_1_net__9_, n_1_net__8_, n_1_net__7_,
         n_1_net__6_, n_1_net__5_, operandA_shift_0_, n_2_net__31_,
         n_2_net__30_, n_2_net__29_, n_2_net__28_, n_2_net__27_, n_2_net__26_,
         n_2_net__25_, n_2_net__24_, n_2_net__23_, n_2_net__22_, n_2_net__21_,
         n_2_net__20_, n_2_net__19_, n_2_net__18_, n_2_net__17_, n_2_net__16_,
         n_2_net__15_, n_2_net__14_, n_2_net__13_, n_2_net__12_, n_2_net__11_,
         n_2_net__10_, n_2_net__9_, n_2_net__8_, n_2_net__7_, n_2_net__6_,
         n_2_net__5_, n_2_net__4_, n_2_net__3_, n_2_net__2_, n_2_net__1_,
         n_2_net__0_, div_sign_ovf, n185, n187, n196, n197, n198, n209, n210,
         n212, n213, n214, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24,
         SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26,
         SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28,
         SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30,
         SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32,
         SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34,
         SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36,
         SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38,
         SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40,
         SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42,
         SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44,
         SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46,
         SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48,
         SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50,
         SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52,
         SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54,
         SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56,
         SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58,
         SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60,
         SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62,
         SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64,
         SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66,
         SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68,
         SYNOPSYS_UNCONNECTED_69, SYNOPSYS_UNCONNECTED_70,
         SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72,
         SYNOPSYS_UNCONNECTED_73, SYNOPSYS_UNCONNECTED_74,
         SYNOPSYS_UNCONNECTED_75, SYNOPSYS_UNCONNECTED_76,
         SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_78,
         SYNOPSYS_UNCONNECTED_79, SYNOPSYS_UNCONNECTED_80,
         SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_82,
         SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_84,
         SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_86,
         SYNOPSYS_UNCONNECTED_87, SYNOPSYS_UNCONNECTED_88,
         SYNOPSYS_UNCONNECTED_89, SYNOPSYS_UNCONNECTED_90,
         SYNOPSYS_UNCONNECTED_91, SYNOPSYS_UNCONNECTED_92,
         SYNOPSYS_UNCONNECTED_93, SYNOPSYS_UNCONNECTED_94,
         SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_96,
         SYNOPSYS_UNCONNECTED_97, SYNOPSYS_UNCONNECTED_98,
         SYNOPSYS_UNCONNECTED_99, SYNOPSYS_UNCONNECTED_100,
         SYNOPSYS_UNCONNECTED_101, SYNOPSYS_UNCONNECTED_102,
         SYNOPSYS_UNCONNECTED_103, SYNOPSYS_UNCONNECTED_104,
         SYNOPSYS_UNCONNECTED_105, SYNOPSYS_UNCONNECTED_106,
         SYNOPSYS_UNCONNECTED_107, SYNOPSYS_UNCONNECTED_108,
         SYNOPSYS_UNCONNECTED_109, SYNOPSYS_UNCONNECTED_110,
         SYNOPSYS_UNCONNECTED_111, SYNOPSYS_UNCONNECTED_112,
         SYNOPSYS_UNCONNECTED_113, SYNOPSYS_UNCONNECTED_114,
         SYNOPSYS_UNCONNECTED_115, SYNOPSYS_UNCONNECTED_116,
         SYNOPSYS_UNCONNECTED_117, SYNOPSYS_UNCONNECTED_118,
         SYNOPSYS_UNCONNECTED_119, SYNOPSYS_UNCONNECTED_120,
         SYNOPSYS_UNCONNECTED_121, SYNOPSYS_UNCONNECTED_122,
         SYNOPSYS_UNCONNECTED_123, SYNOPSYS_UNCONNECTED_124,
         SYNOPSYS_UNCONNECTED_125, SYNOPSYS_UNCONNECTED_126,
         SYNOPSYS_UNCONNECTED_127, SYNOPSYS_UNCONNECTED_128,
         \ctrl/SYNOPSYS_UNCONNECTED_2 , \ctrl/SYNOPSYS_UNCONNECTED_1 ,
         \ctrl/n22 , \ctrl/n21 , \ctrl/n20 , \ctrl/n19 , \ctrl/n18 ,
         \ctrl/n17 , \ctrl/n15 , \ctrl/n14 , \ctrl/n13 , \ctrl/n12 ,
         \ctrl/n11 , \ctrl/n10 , \ctrl/n9 , \ctrl/n8 , \ctrl/n7 ,
         \ctrl/n_3_net_ , \ctrl/op_div_int , \ctrl/mult_ready ,
         \ctrl/op_mult_int , \ctrl/decoded_seq[1] , \ctrl/decoded_seq[2] ,
         \ctrl/decoded_seq[3] , \ctrl/decoded_seq[4] , \ctrl/decoded_seq[5] ,
         \ctrl/decoded_seq[6] , \ctrl/decoder/n11 , \ctrl/decoder/n10 ,
         \ctrl/decoder/n9 , \ctrl/decoder/n8 , \ctrl/decoder/n7 ,
         \ctrl/decoder/n6 , \ctrl/decoder/n5 , \ctrl/decoder/n4 ,
         \ctrl/decoder/n3 , \ctrl/decoder/n2 , \ctrl/decoder/n1 ,
         \ctrl/counter/n1 , \ctrl/counter/w7 , \ctrl/counter/w6 ,
         \ctrl/counter/w5 , \ctrl/counter/w4 , \ctrl/counter/w3 ,
         \ctrl/counter/w2 , \ctrl/counter/w1 , \ctrl/counter/tff_0/d ,
         \ctrl/counter/tff_0/data , \ctrl/counter/tff_0/dffe/n7 ,
         \ctrl/counter/tff_0/dffe/n6 , \ctrl/counter/tff_0/dffe/n5 ,
         \ctrl/counter/tff_0/dffe/n1 , \ctrl/counter/tff_1/d ,
         \ctrl/counter/tff_1/data , \ctrl/counter/tff_1/dffe/n7 ,
         \ctrl/counter/tff_1/dffe/n6 , \ctrl/counter/tff_1/dffe/n5 ,
         \ctrl/counter/tff_1/dffe/n1 , \ctrl/counter/tff_2/d ,
         \ctrl/counter/tff_2/data , \ctrl/counter/tff_2/dffe/n7 ,
         \ctrl/counter/tff_2/dffe/n6 , \ctrl/counter/tff_2/dffe/n5 ,
         \ctrl/counter/tff_2/dffe/n1 , \ctrl/counter/tff_3/d ,
         \ctrl/counter/tff_3/data , \ctrl/counter/tff_3/dffe/n7 ,
         \ctrl/counter/tff_3/dffe/n6 , \ctrl/counter/tff_3/dffe/n5 ,
         \ctrl/counter/tff_3/dffe/n1 , \ctrl/counter/tff_4/d ,
         \ctrl/counter/tff_4/dffe/n7 , \ctrl/counter/tff_4/dffe/n6 ,
         \ctrl/counter/tff_4/dffe/n5 , \ctrl/counter/tff_4/dffe/n1 ,
         \ctrl/counter/tff_5/data_not , \ctrl/counter/tff_5/d ,
         \ctrl/counter/tff_5/dffe/n7 , \ctrl/counter/tff_5/dffe/n6 ,
         \ctrl/counter/tff_5/dffe/n5 , \ctrl/counter/tff_5/dffe/n1 ,
         \ctrl/counter/output16_dff/n7 , \ctrl/counter/output16_dff/n6 ,
         \ctrl/counter/output16_dff/n5 , \ctrl/counter/output16_dff/n1 ,
         \ctrl/counter/output32_dff/n7 , \ctrl/counter/output32_dff/n6 ,
         \ctrl/counter/output32_dff/n5 , \ctrl/counter/output32_dff/n1 ,
         \ctrl/cur_mult/n4 , \ctrl/cur_mult/n3 , \ctrl/cur_mult/n2 ,
         \ctrl/cur_mult/n1 , \ctrl/cur_div/n7 , \ctrl/cur_div/n6 ,
         \ctrl/cur_div/n5 , \ctrl/cur_div/n1 , \add_sub_mux/n76 ,
         \add_sub_mux/n75 , \add_sub_mux/n74 , \add_sub_mux/n73 ,
         \add_sub_mux/n72 , \add_sub_mux/n71 , \add_sub_mux/n70 ,
         \add_sub_mux/n69 , \add_sub_mux/n68 , \add_sub_mux/n67 ,
         \add_sub_mux/n66 , \add_sub_mux/n33 , \add_sub_mux/n65 ,
         \add_sub_mux/n64 , \add_sub_mux/n63 , \add_sub_mux/n62 ,
         \add_sub_mux/n61 , \add_sub_mux/n60 , \add_sub_mux/n59 ,
         \add_sub_mux/n58 , \add_sub_mux/n57 , \add_sub_mux/n56 ,
         \add_sub_mux/n55 , \add_sub_mux/n54 , \add_sub_mux/n53 ,
         \add_sub_mux/n52 , \add_sub_mux/n51 , \add_sub_mux/n50 ,
         \add_sub_mux/n49 , \add_sub_mux/n48 , \add_sub_mux/n47 ,
         \add_sub_mux/n46 , \add_sub_mux/n45 , \add_sub_mux/n44 ,
         \add_sub_mux/n43 , \add_sub_mux/n42 , \add_sub_mux/n41 ,
         \add_sub_mux/n40 , \add_sub_mux/n39 , \add_sub_mux/n38 ,
         \add_sub_mux/n37 , \add_sub_mux/n36 , \add_sub_mux/n35 ,
         \add_sub_mux/n34 , \shift_booth_mux/n101 , \shift_booth_mux/n100 ,
         \shift_booth_mux/n99 , \shift_booth_mux/n98 , \shift_booth_mux/n97 ,
         \shift_booth_mux/n96 , \shift_booth_mux/n95 , \shift_booth_mux/n94 ,
         \shift_booth_mux/n93 , \shift_booth_mux/n92 , \shift_booth_mux/n91 ,
         \shift_booth_mux/n90 , \shift_booth_mux/n89 , \shift_booth_mux/n88 ,
         \shift_booth_mux/n87 , \shift_booth_mux/n86 , \shift_booth_mux/n85 ,
         \shift_booth_mux/n84 , \shift_booth_mux/n83 , \shift_booth_mux/n82 ,
         \shift_booth_mux/n81 , \shift_booth_mux/n80 , \shift_booth_mux/n79 ,
         \shift_booth_mux/n78 , \shift_booth_mux/n77 , \shift_booth_mux/n76 ,
         \shift_booth_mux/n75 , \shift_booth_mux/n74 , \shift_booth_mux/n73 ,
         \shift_booth_mux/n72 , \shift_booth_mux/n71 , \shift_booth_mux/n70 ,
         \shift_booth_mux/n69 , \shift_booth_mux/n68 , \shift_booth_mux/n67 ,
         \shift_booth_mux/n66 , \shift_booth_mux/n65 , \shift_booth_mux/n54 ,
         \shift_booth_mux/n43 , \shift_booth_mux/n40 , \shift_booth_mux/n33 ,
         \nop_mux/n100 , \nop_mux/n99 , \nop_mux/n98 , \nop_mux/n97 ,
         \nop_mux/n96 , \nop_mux/n95 , \nop_mux/n94 , \nop_mux/n93 ,
         \nop_mux/n92 , \nop_mux/n91 , \nop_mux/n90 , \nop_mux/n89 ,
         \nop_mux/n88 , \nop_mux/n87 , \nop_mux/n86 , \nop_mux/n85 ,
         \nop_mux/n84 , \nop_mux/n83 , \nop_mux/n82 , \nop_mux/n81 ,
         \nop_mux/n80 , \nop_mux/n79 , \nop_mux/n78 , \nop_mux/n77 ,
         \nop_mux/n76 , \nop_mux/n75 , \nop_mux/n74 , \nop_mux/n73 ,
         \nop_mux/n72 , \nop_mux/n71 , \nop_mux/n70 , \nop_mux/n69 ,
         \nop_mux/n68 , \nop_mux/n67 , \nop_mux/n66 , \nop_mux/n65 ,
         \nop_mux/n54 , \nop_mux/n43 , \nop_mux/n33 , \adder/n18 , \adder/n17 ,
         \adder/n16 , \adder/n15 , \adder/n14 , \adder/n13 , \adder/n12 ,
         \adder/n11 , \adder/n10 , \adder/g2 , \adder/p2 , \adder/g1 ,
         \adder/p1 , \adder/g0 , \adder/p0 , \adder/overflow ,
         \adder/adder1/n86 , \adder/adder1/n85 , \adder/adder1/n84 ,
         \adder/adder1/n83 , \adder/adder1/n82 , \adder/adder1/n81 ,
         \adder/adder1/n80 , \adder/adder1/n79 , \adder/adder1/n78 ,
         \adder/adder1/n77 , \adder/adder1/n75 , \adder/adder1/n74 ,
         \adder/adder1/n72 , \adder/adder1/n71 , \adder/adder1/n70 ,
         \adder/adder1/n69 , \adder/adder1/n68 , \adder/adder1/n64 ,
         \adder/adder1/n63 , \adder/adder1/n62 , \adder/adder1/n60 ,
         \adder/adder1/n49 , \adder/adder1/n59 , \adder/adder1/n58 ,
         \adder/adder1/n57 , \adder/adder1/n55 , \adder/adder1/n54 ,
         \adder/adder1/n53 , \adder/adder1/n52 , \adder/adder1/n51 ,
         \adder/adder1/n50 , \adder/adder1/n48 , \adder/adder1/n47 ,
         \adder/adder1/n46 , \adder/adder1/n45 , \adder/adder1/n44 ,
         \adder/adder1/n43 , \adder/adder1/n42 , \adder/adder1/n41 ,
         \adder/adder1/n40 , \adder/adder1/n39 , \adder/adder1/n38 ,
         \adder/adder1/n37 , \adder/adder1/n36 , \adder/adder1/n35 ,
         \adder/adder1/n34 , \adder/adder1/n33 , \adder/adder1/n32 ,
         \adder/adder1/n31 , \adder/adder1/n30 , \adder/adder1/n29 ,
         \adder/adder1/n28 , \adder/adder1/n27 , \adder/adder1/n26 ,
         \adder/adder1/n17 , \adder/adder1/n15 , \adder/adder1/n14 ,
         \adder/adder1/n13 , \adder/adder1/n87 , \adder/adder1/overflow ,
         \adder/adder1/n88 , \adder/adder2/n110 , \adder/adder2/n109 ,
         \adder/adder2/n107 , \adder/adder2/n106 , \adder/adder2/n105 ,
         \adder/adder2/n104 , \adder/adder2/n103 , \adder/adder2/n102 ,
         \adder/adder2/n101 , \adder/adder2/n100 , \adder/adder2/n99 ,
         \adder/adder2/n98 , \adder/adder2/n97 , \adder/adder2/n96 ,
         \adder/adder2/n95 , \adder/adder2/n94 , \adder/adder2/n93 ,
         \adder/adder2/n92 , \adder/adder2/n91 , \adder/adder2/n90 ,
         \adder/adder2/n89 , \adder/adder2/n88 , \adder/adder2/n87 ,
         \adder/adder2/n86 , \adder/adder2/n85 , \adder/adder2/n84 ,
         \adder/adder2/n83 , \adder/adder2/n82 , \adder/adder2/n81 ,
         \adder/adder2/n80 , \adder/adder2/n79 , \adder/adder2/n78 ,
         \adder/adder2/n77 , \adder/adder2/n76 , \adder/adder2/n75 ,
         \adder/adder2/n74 , \adder/adder2/n73 , \adder/adder2/n72 ,
         \adder/adder2/n71 , \adder/adder2/n70 , \adder/adder2/n69 ,
         \adder/adder2/n68 , \adder/adder2/n67 , \adder/adder2/n66 ,
         \adder/adder2/n65 , \adder/adder2/n64 , \adder/adder2/n63 ,
         \adder/adder2/n62 , \adder/adder2/n61 , \adder/adder2/n60 ,
         \adder/adder2/n56 , \adder/adder2/overflow , \adder/adder3/n110 ,
         \adder/adder3/n109 , \adder/adder3/n107 , \adder/adder3/n106 ,
         \adder/adder3/n105 , \adder/adder3/n104 , \adder/adder3/n103 ,
         \adder/adder3/n102 , \adder/adder3/n101 , \adder/adder3/n100 ,
         \adder/adder3/n99 , \adder/adder3/n98 , \adder/adder3/n97 ,
         \adder/adder3/n96 , \adder/adder3/n95 , \adder/adder3/n94 ,
         \adder/adder3/n93 , \adder/adder3/n92 , \adder/adder3/n91 ,
         \adder/adder3/n90 , \adder/adder3/n89 , \adder/adder3/n88 ,
         \adder/adder3/n87 , \adder/adder3/n86 , \adder/adder3/n85 ,
         \adder/adder3/n84 , \adder/adder3/n83 , \adder/adder3/n82 ,
         \adder/adder3/n81 , \adder/adder3/n80 , \adder/adder3/n79 ,
         \adder/adder3/n78 , \adder/adder3/n77 , \adder/adder3/n76 ,
         \adder/adder3/n75 , \adder/adder3/n74 , \adder/adder3/n73 ,
         \adder/adder3/n72 , \adder/adder3/n71 , \adder/adder3/n70 ,
         \adder/adder3/n69 , \adder/adder3/n68 , \adder/adder3/n67 ,
         \adder/adder3/n66 , \adder/adder3/n65 , \adder/adder3/n64 ,
         \adder/adder3/n63 , \adder/adder3/n62 , \adder/adder3/n61 ,
         \adder/adder3/n60 , \adder/adder3/n56 , \adder/adder3/overflow ,
         \adder/adder4/n111 , \adder/adder4/n110 , \adder/adder4/n109 ,
         \adder/adder4/n108 , \adder/adder4/n107 , \adder/adder4/n106 ,
         \adder/adder4/n105 , \adder/adder4/n104 , \adder/adder4/n103 ,
         \adder/adder4/n102 , \adder/adder4/n101 , \adder/adder4/n100 ,
         \adder/adder4/n99 , \adder/adder4/n98 , \adder/adder4/n97 ,
         \adder/adder4/n96 , \adder/adder4/n95 , \adder/adder4/n94 ,
         \adder/adder4/n93 , \adder/adder4/n92 , \adder/adder4/n91 ,
         \adder/adder4/n90 , \adder/adder4/n89 , \adder/adder4/n88 ,
         \adder/adder4/n87 , \adder/adder4/n86 , \adder/adder4/n85 ,
         \adder/adder4/n84 , \adder/adder4/n83 , \adder/adder4/n82 ,
         \adder/adder4/n81 , \adder/adder4/n80 , \adder/adder4/n79 ,
         \adder/adder4/n78 , \adder/adder4/n77 , \adder/adder4/n76 ,
         \adder/adder4/n75 , \adder/adder4/n74 , \adder/adder4/n73 ,
         \adder/adder4/n72 , \adder/adder4/n71 , \adder/adder4/n70 ,
         \adder/adder4/n69 , \adder/adder4/n68 , \adder/adder4/n67 ,
         \adder/adder4/n66 , \adder/adder4/n65 , \adder/adder4/n64 ,
         \adder/adder4/n63 , \adder/adder4/n62 , \adder/adder4/n61 ,
         \adder/adder4/n60 , \adder/adder4/gen , \adder/adder4/prop ,
         \adder_sign/n17 , \adder_sign/n16 , \adder_sign/n15 ,
         \adder_sign/n14 , \adder_sign/n13 , \adder_sign/n12 ,
         \adder_sign/n11 , \adder_sign/n10 , \adder_sign/g2 , \adder_sign/p2 ,
         \adder_sign/g1 , \adder_sign/p1 , \adder_sign/g0 , \adder_sign/p0 ,
         \adder_sign/adder1/n104 , \adder_sign/adder1/n103 ,
         \adder_sign/adder1/n101 , \adder_sign/adder1/n100 ,
         \adder_sign/adder1/n99 , \adder_sign/adder1/n98 ,
         \adder_sign/adder1/n97 , \adder_sign/adder1/n96 ,
         \adder_sign/adder1/n95 , \adder_sign/adder1/n94 ,
         \adder_sign/adder1/n93 , \adder_sign/adder1/n92 ,
         \adder_sign/adder1/n91 , \adder_sign/adder1/n90 ,
         \adder_sign/adder1/n89 , \adder_sign/adder1/n88 ,
         \adder_sign/adder1/n87 , \adder_sign/adder1/n86 ,
         \adder_sign/adder1/n85 , \adder_sign/adder1/n84 ,
         \adder_sign/adder1/n83 , \adder_sign/adder1/n82 ,
         \adder_sign/adder1/n81 , \adder_sign/adder1/n80 ,
         \adder_sign/adder1/n79 , \adder_sign/adder1/n78 ,
         \adder_sign/adder1/n77 , \adder_sign/adder1/n76 ,
         \adder_sign/adder1/n75 , \adder_sign/adder1/n74 ,
         \adder_sign/adder1/n73 , \adder_sign/adder1/n72 ,
         \adder_sign/adder1/n71 , \adder_sign/adder1/n70 ,
         \adder_sign/adder1/n69 , \adder_sign/adder1/n68 ,
         \adder_sign/adder1/n67 , \adder_sign/adder1/n66 ,
         \adder_sign/adder1/n65 , \adder_sign/adder1/n64 ,
         \adder_sign/adder1/n63 , \adder_sign/adder1/n62 ,
         \adder_sign/adder1/n61 , \adder_sign/adder1/n60 ,
         \adder_sign/adder1/overflow , \adder_sign/adder2/n105 ,
         \adder_sign/adder2/n104 , \adder_sign/adder2/n103 ,
         \adder_sign/adder2/n102 , \adder_sign/adder2/n101 ,
         \adder_sign/adder2/n100 , \adder_sign/adder2/n99 ,
         \adder_sign/adder2/n98 , \adder_sign/adder2/n97 ,
         \adder_sign/adder2/n96 , \adder_sign/adder2/n95 ,
         \adder_sign/adder2/n94 , \adder_sign/adder2/n93 ,
         \adder_sign/adder2/n92 , \adder_sign/adder2/n91 ,
         \adder_sign/adder2/n90 , \adder_sign/adder2/n89 ,
         \adder_sign/adder2/n88 , \adder_sign/adder2/n87 ,
         \adder_sign/adder2/n86 , \adder_sign/adder2/n85 ,
         \adder_sign/adder2/n84 , \adder_sign/adder2/n83 ,
         \adder_sign/adder2/n82 , \adder_sign/adder2/n81 ,
         \adder_sign/adder2/n80 , \adder_sign/adder2/n79 ,
         \adder_sign/adder2/n78 , \adder_sign/adder2/n77 ,
         \adder_sign/adder2/n76 , \adder_sign/adder2/n75 ,
         \adder_sign/adder2/n74 , \adder_sign/adder2/n73 ,
         \adder_sign/adder2/n72 , \adder_sign/adder2/n71 ,
         \adder_sign/adder2/n70 , \adder_sign/adder2/n69 ,
         \adder_sign/adder2/n68 , \adder_sign/adder2/n67 ,
         \adder_sign/adder2/n66 , \adder_sign/adder2/n65 ,
         \adder_sign/adder2/n64 , \adder_sign/adder2/n63 ,
         \adder_sign/adder2/n62 , \adder_sign/adder2/n61 ,
         \adder_sign/adder2/n60 , \adder_sign/adder2/overflow ,
         \adder_sign/adder3/n104 , \adder_sign/adder3/n103 ,
         \adder_sign/adder3/n102 , \adder_sign/adder3/n101 ,
         \adder_sign/adder3/n100 , \adder_sign/adder3/n99 ,
         \adder_sign/adder3/n98 , \adder_sign/adder3/n97 ,
         \adder_sign/adder3/n96 , \adder_sign/adder3/n95 ,
         \adder_sign/adder3/n94 , \adder_sign/adder3/n93 ,
         \adder_sign/adder3/n92 , \adder_sign/adder3/n91 ,
         \adder_sign/adder3/n90 , \adder_sign/adder3/n89 ,
         \adder_sign/adder3/n88 , \adder_sign/adder3/n87 ,
         \adder_sign/adder3/n86 , \adder_sign/adder3/n85 ,
         \adder_sign/adder3/n84 , \adder_sign/adder3/n83 ,
         \adder_sign/adder3/n82 , \adder_sign/adder3/n81 ,
         \adder_sign/adder3/n80 , \adder_sign/adder3/n79 ,
         \adder_sign/adder3/n78 , \adder_sign/adder3/n77 ,
         \adder_sign/adder3/n76 , \adder_sign/adder3/n75 ,
         \adder_sign/adder3/n74 , \adder_sign/adder3/n73 ,
         \adder_sign/adder3/n72 , \adder_sign/adder3/n71 ,
         \adder_sign/adder3/n70 , \adder_sign/adder3/n69 ,
         \adder_sign/adder3/n68 , \adder_sign/adder3/n67 ,
         \adder_sign/adder3/n66 , \adder_sign/adder3/n65 ,
         \adder_sign/adder3/n64 , \adder_sign/adder3/n63 ,
         \adder_sign/adder3/n62 , \adder_sign/adder3/n61 ,
         \adder_sign/adder3/n60 , \adder_sign/adder3/overflow ,
         \adder_sign/adder4/n103 , \adder_sign/adder4/n102 ,
         \adder_sign/adder4/n101 , \adder_sign/adder4/n100 ,
         \adder_sign/adder4/n99 , \adder_sign/adder4/n98 ,
         \adder_sign/adder4/n97 , \adder_sign/adder4/n96 ,
         \adder_sign/adder4/n95 , \adder_sign/adder4/n94 ,
         \adder_sign/adder4/n93 , \adder_sign/adder4/n92 ,
         \adder_sign/adder4/n91 , \adder_sign/adder4/n90 ,
         \adder_sign/adder4/n89 , \adder_sign/adder4/n88 ,
         \adder_sign/adder4/n87 , \adder_sign/adder4/n86 ,
         \adder_sign/adder4/n85 , \adder_sign/adder4/n84 ,
         \adder_sign/adder4/n83 , \adder_sign/adder4/n82 ,
         \adder_sign/adder4/n81 , \adder_sign/adder4/n80 ,
         \adder_sign/adder4/n79 , \adder_sign/adder4/n78 ,
         \adder_sign/adder4/n77 , \adder_sign/adder4/n76 ,
         \adder_sign/adder4/n75 , \adder_sign/adder4/n74 ,
         \adder_sign/adder4/n73 , \adder_sign/adder4/n72 ,
         \adder_sign/adder4/n71 , \adder_sign/adder4/n70 ,
         \adder_sign/adder4/n69 , \adder_sign/adder4/n68 ,
         \adder_sign/adder4/n67 , \adder_sign/adder4/n66 ,
         \adder_sign/adder4/n65 , \adder_sign/adder4/n64 ,
         \adder_sign/adder4/n63 , \adder_sign/adder4/n62 ,
         \adder_sign/adder4/n61 , \adder_sign/adder4/n60 ,
         \adder_sign/adder4/gen , \adder_sign/adder4/prop , \product_reg/n7 ,
         \product_reg/n6 , \product_reg/n5 , \product_reg/n4 ,
         \product_reg/n3 , \product_reg/n2 , \product_reg/n1 ,
         \product_reg/memory_0__dff/n7 , \product_reg/memory_0__dff/n6 ,
         \product_reg/memory_0__dff/n5 , \product_reg/memory_0__dff/n1 ,
         \product_reg/memory_1__dff/n10 , \product_reg/memory_1__dff/n9 ,
         \product_reg/memory_1__dff/n8 , \product_reg/memory_1__dff/n6 ,
         \product_reg/memory_1__dff/n5 , \product_reg/memory_1__dff/n1 ,
         \product_reg/memory_2__dff/n10 , \product_reg/memory_2__dff/n9 ,
         \product_reg/memory_2__dff/n7 , \product_reg/memory_2__dff/n4 ,
         \product_reg/memory_2__dff/n1 , \product_reg/memory_3__dff/n7 ,
         \product_reg/memory_3__dff/n6 , \product_reg/memory_3__dff/n5 ,
         \product_reg/memory_3__dff/n1 , \product_reg/memory_4__dff/n7 ,
         \product_reg/memory_4__dff/n6 , \product_reg/memory_4__dff/n5 ,
         \product_reg/memory_4__dff/n1 , \product_reg/memory_5__dff/n7 ,
         \product_reg/memory_5__dff/n6 , \product_reg/memory_5__dff/n5 ,
         \product_reg/memory_5__dff/n1 , \product_reg/memory_6__dff/n7 ,
         \product_reg/memory_6__dff/n6 , \product_reg/memory_6__dff/n5 ,
         \product_reg/memory_6__dff/n1 , \product_reg/memory_7__dff/n7 ,
         \product_reg/memory_7__dff/n6 , \product_reg/memory_7__dff/n5 ,
         \product_reg/memory_7__dff/n1 , \product_reg/memory_8__dff/n7 ,
         \product_reg/memory_8__dff/n6 , \product_reg/memory_8__dff/n5 ,
         \product_reg/memory_8__dff/n1 , \product_reg/memory_9__dff/n7 ,
         \product_reg/memory_9__dff/n6 , \product_reg/memory_9__dff/n5 ,
         \product_reg/memory_9__dff/n1 , \product_reg/memory_10__dff/n7 ,
         \product_reg/memory_10__dff/n6 , \product_reg/memory_10__dff/n5 ,
         \product_reg/memory_10__dff/n1 , \product_reg/memory_11__dff/n7 ,
         \product_reg/memory_11__dff/n6 , \product_reg/memory_11__dff/n5 ,
         \product_reg/memory_11__dff/n1 , \product_reg/memory_12__dff/n7 ,
         \product_reg/memory_12__dff/n6 , \product_reg/memory_12__dff/n5 ,
         \product_reg/memory_12__dff/n1 , \product_reg/memory_13__dff/n7 ,
         \product_reg/memory_13__dff/n6 , \product_reg/memory_13__dff/n5 ,
         \product_reg/memory_13__dff/n1 , \product_reg/memory_14__dff/n7 ,
         \product_reg/memory_14__dff/n6 , \product_reg/memory_14__dff/n5 ,
         \product_reg/memory_14__dff/n1 , \product_reg/memory_15__dff/n7 ,
         \product_reg/memory_15__dff/n6 , \product_reg/memory_15__dff/n5 ,
         \product_reg/memory_15__dff/n1 , \product_reg/memory_16__dff/n7 ,
         \product_reg/memory_16__dff/n6 , \product_reg/memory_16__dff/n5 ,
         \product_reg/memory_16__dff/n1 , \product_reg/memory_17__dff/n7 ,
         \product_reg/memory_17__dff/n6 , \product_reg/memory_17__dff/n5 ,
         \product_reg/memory_17__dff/n1 , \product_reg/memory_18__dff/n7 ,
         \product_reg/memory_18__dff/n6 , \product_reg/memory_18__dff/n5 ,
         \product_reg/memory_18__dff/n1 , \product_reg/memory_19__dff/n7 ,
         \product_reg/memory_19__dff/n6 , \product_reg/memory_19__dff/n5 ,
         \product_reg/memory_19__dff/n1 , \product_reg/memory_20__dff/n7 ,
         \product_reg/memory_20__dff/n6 , \product_reg/memory_20__dff/n5 ,
         \product_reg/memory_20__dff/n1 , \product_reg/memory_21__dff/n7 ,
         \product_reg/memory_21__dff/n6 , \product_reg/memory_21__dff/n5 ,
         \product_reg/memory_21__dff/n1 , \product_reg/memory_22__dff/n7 ,
         \product_reg/memory_22__dff/n6 , \product_reg/memory_22__dff/n5 ,
         \product_reg/memory_22__dff/n1 , \product_reg/memory_23__dff/n7 ,
         \product_reg/memory_23__dff/n6 , \product_reg/memory_23__dff/n5 ,
         \product_reg/memory_23__dff/n1 , \product_reg/memory_24__dff/n7 ,
         \product_reg/memory_24__dff/n6 , \product_reg/memory_24__dff/n5 ,
         \product_reg/memory_24__dff/n1 , \product_reg/memory_25__dff/n7 ,
         \product_reg/memory_25__dff/n6 , \product_reg/memory_25__dff/n5 ,
         \product_reg/memory_25__dff/n1 , \product_reg/memory_26__dff/n7 ,
         \product_reg/memory_26__dff/n6 , \product_reg/memory_26__dff/n5 ,
         \product_reg/memory_26__dff/n1 , \product_reg/memory_27__dff/n7 ,
         \product_reg/memory_27__dff/n6 , \product_reg/memory_27__dff/n5 ,
         \product_reg/memory_27__dff/n1 , \product_reg/memory_28__dff/n7 ,
         \product_reg/memory_28__dff/n6 , \product_reg/memory_28__dff/n5 ,
         \product_reg/memory_28__dff/n1 , \product_reg/memory_29__dff/n7 ,
         \product_reg/memory_29__dff/n6 , \product_reg/memory_29__dff/n5 ,
         \product_reg/memory_29__dff/n1 , \product_reg/memory_30__dff/n7 ,
         \product_reg/memory_30__dff/n6 , \product_reg/memory_30__dff/n5 ,
         \product_reg/memory_30__dff/n1 , \product_reg/memory_31__dff/n7 ,
         \product_reg/memory_31__dff/n6 , \product_reg/memory_31__dff/n5 ,
         \product_reg/memory_31__dff/n1 , \product_reg/memory_32__dff/n3 ,
         \product_reg/memory_32__dff/n1 , \product_reg/memory_33__dff/n7 ,
         \product_reg/memory_33__dff/n6 , \product_reg/memory_33__dff/n5 ,
         \product_reg/memory_33__dff/n1 , \product_reg/memory_34__dff/n7 ,
         \product_reg/memory_34__dff/n6 , \product_reg/memory_34__dff/n5 ,
         \product_reg/memory_34__dff/n1 , \product_reg/memory_35__dff/n7 ,
         \product_reg/memory_35__dff/n6 , \product_reg/memory_35__dff/n5 ,
         \product_reg/memory_35__dff/n1 , \product_reg/memory_36__dff/n7 ,
         \product_reg/memory_36__dff/n6 , \product_reg/memory_36__dff/n5 ,
         \product_reg/memory_36__dff/n1 , \product_reg/memory_37__dff/n7 ,
         \product_reg/memory_37__dff/n6 , \product_reg/memory_37__dff/n5 ,
         \product_reg/memory_37__dff/n1 , \product_reg/memory_38__dff/n7 ,
         \product_reg/memory_38__dff/n6 , \product_reg/memory_38__dff/n5 ,
         \product_reg/memory_38__dff/n1 , \product_reg/memory_39__dff/n7 ,
         \product_reg/memory_39__dff/n6 , \product_reg/memory_39__dff/n5 ,
         \product_reg/memory_39__dff/n1 , \product_reg/memory_40__dff/n7 ,
         \product_reg/memory_40__dff/n6 , \product_reg/memory_40__dff/n5 ,
         \product_reg/memory_40__dff/n1 , \product_reg/memory_41__dff/n7 ,
         \product_reg/memory_41__dff/n6 , \product_reg/memory_41__dff/n5 ,
         \product_reg/memory_41__dff/n1 , \product_reg/memory_42__dff/n7 ,
         \product_reg/memory_42__dff/n6 , \product_reg/memory_42__dff/n5 ,
         \product_reg/memory_42__dff/n1 , \product_reg/memory_43__dff/n7 ,
         \product_reg/memory_43__dff/n6 , \product_reg/memory_43__dff/n5 ,
         \product_reg/memory_43__dff/n1 , \product_reg/memory_44__dff/n7 ,
         \product_reg/memory_44__dff/n6 , \product_reg/memory_44__dff/n5 ,
         \product_reg/memory_44__dff/n1 , \product_reg/memory_45__dff/n7 ,
         \product_reg/memory_45__dff/n6 , \product_reg/memory_45__dff/n5 ,
         \product_reg/memory_45__dff/n1 , \product_reg/memory_46__dff/n7 ,
         \product_reg/memory_46__dff/n6 , \product_reg/memory_46__dff/n5 ,
         \product_reg/memory_46__dff/n1 , \product_reg/memory_47__dff/n7 ,
         \product_reg/memory_47__dff/n6 , \product_reg/memory_47__dff/n5 ,
         \product_reg/memory_47__dff/n1 , \product_reg/memory_48__dff/n7 ,
         \product_reg/memory_48__dff/n6 , \product_reg/memory_48__dff/n5 ,
         \product_reg/memory_48__dff/n1 , \product_reg/memory_49__dff/n7 ,
         \product_reg/memory_49__dff/n6 , \product_reg/memory_49__dff/n5 ,
         \product_reg/memory_49__dff/n1 , \product_reg/memory_50__dff/n7 ,
         \product_reg/memory_50__dff/n6 , \product_reg/memory_50__dff/n5 ,
         \product_reg/memory_50__dff/n1 , \product_reg/memory_51__dff/n7 ,
         \product_reg/memory_51__dff/n6 , \product_reg/memory_51__dff/n5 ,
         \product_reg/memory_51__dff/n1 , \product_reg/memory_52__dff/n7 ,
         \product_reg/memory_52__dff/n6 , \product_reg/memory_52__dff/n5 ,
         \product_reg/memory_52__dff/n1 , \product_reg/memory_53__dff/n7 ,
         \product_reg/memory_53__dff/n6 , \product_reg/memory_53__dff/n5 ,
         \product_reg/memory_53__dff/n1 , \product_reg/memory_54__dff/n7 ,
         \product_reg/memory_54__dff/n6 , \product_reg/memory_54__dff/n5 ,
         \product_reg/memory_54__dff/n1 , \product_reg/memory_55__dff/n7 ,
         \product_reg/memory_55__dff/n6 , \product_reg/memory_55__dff/n5 ,
         \product_reg/memory_55__dff/n1 , \product_reg/memory_56__dff/n7 ,
         \product_reg/memory_56__dff/n6 , \product_reg/memory_56__dff/n5 ,
         \product_reg/memory_56__dff/n1 , \product_reg/memory_57__dff/n7 ,
         \product_reg/memory_57__dff/n6 , \product_reg/memory_57__dff/n5 ,
         \product_reg/memory_57__dff/n1 , \product_reg/memory_58__dff/n7 ,
         \product_reg/memory_58__dff/n6 , \product_reg/memory_58__dff/n5 ,
         \product_reg/memory_58__dff/n1 , \product_reg/memory_59__dff/n7 ,
         \product_reg/memory_59__dff/n6 , \product_reg/memory_59__dff/n5 ,
         \product_reg/memory_59__dff/n1 , \product_reg/memory_60__dff/n7 ,
         \product_reg/memory_60__dff/n6 , \product_reg/memory_60__dff/n5 ,
         \product_reg/memory_60__dff/n1 , \product_reg/memory_61__dff/n7 ,
         \product_reg/memory_61__dff/n6 , \product_reg/memory_61__dff/n5 ,
         \product_reg/memory_61__dff/n1 , \product_reg/memory_62__dff/n7 ,
         \product_reg/memory_62__dff/n6 , \product_reg/memory_62__dff/n5 ,
         \product_reg/memory_62__dff/n1 , \product_reg/memory_63__dff/n8 ,
         \product_reg/memory_63__dff/n7 , \product_reg/memory_63__dff/n6 ,
         \product_reg/memory_63__dff/n5 , \product_reg/memory_63__dff/n1 ,
         \product_reg/memory_64__dff/n7 , \product_reg/memory_64__dff/n6 ,
         \product_reg/memory_64__dff/n5 , \product_reg/memory_64__dff/n1 ;
  wire   [64:0] product_out;
  wire   [31:0] data_operandA_not;
  wire   [31:0] operandA;
  wire   [31:0] operandA_resolved;
  wire   [31:0] alu_operand;
  wire   [31:0] adder_out;
  wire   [31:0] sign_fixed;
  wire   [64:0] product_in;

  NAND3_X1 U708 ( .A1(n508), .A2(n507), .A3(n509), .ZN(n535) );
  NAND3_X1 U709 ( .A1(n438), .A2(n439), .A3(n437), .ZN(n545) );
  NAND3_X1 U710 ( .A1(product_out[33]), .A2(product_out[32]), .A3(
        product_out[34]), .ZN(n555) );
  XOR2_X1 U711 ( .A(data_operandB[31]), .B(n681), .Z(n522) );
  TBUF_X1 product_in_tri_62_ ( .A(adder_out[31]), .EN(n630), .Z(product_in[62]) );
  TBUF_X1 product_in_tri4_62_ ( .A(adder_out[29]), .EN(n340), .Z(
        product_in[62]) );
  TBUF_X1 product_in_tri3_62_ ( .A(1'b0), .EN(n677), .Z(product_in[62]) );
  TBUF_X1 product_in_tri2_62_ ( .A(1'b0), .EN(n635), .Z(product_in[62]) );
  TBUF_X1 product_in_tri_64_ ( .A(n625), .EN(n630), .Z(product_in[64]) );
  TBUF_X1 product_in_tri4_3_ ( .A(n624), .EN(n340), .Z(product_in[3]) );
  TBUF_X1 product_in_tri_0_ ( .A(n624), .EN(n654), .Z(product_in[0]) );
  TBUF_X1 product_in_tri4_2_ ( .A(n619), .EN(n340), .Z(product_in[2]) );
  TBUF_X1 product_in_tri4_33_ ( .A(adder_out[0]), .EN(n640), .Z(product_in[33]) );
  TBUF_X1 product_in_tri_31_ ( .A(adder_out[0]), .EN(n618), .Z(product_in[31])
         );
  TBUF_X1 product_in_tri_63_ ( .A(n185), .EN(n618), .Z(product_in[63]) );
  TBUF_X1 product_in_tri2_63_ ( .A(1'b0), .EN(n636), .Z(product_in[63]) );
  TBUF_X1 product_in_tri3_63_ ( .A(1'b0), .EN(n679), .Z(product_in[63]) );
  TBUF_X1 product_in_tri4_63_ ( .A(adder_out[30]), .EN(n340), .Z(
        product_in[63]) );
  TBUF_X1 product_in_tri_33_ ( .A(adder_out[2]), .EN(n618), .Z(product_in[33])
         );
  TBUF_X1 product_in_tri_32_ ( .A(adder_out[1]), .EN(n618), .Z(product_in[32])
         );
  TBUF_X1 product_in_tri_34_ ( .A(adder_out[3]), .EN(n618), .Z(product_in[34])
         );
  TBUF_X1 product_in_tri4_7_ ( .A(product_out[6]), .EN(n340), .Z(product_in[7]) );
  TBUF_X1 product_in_tri4_8_ ( .A(product_out[7]), .EN(n340), .Z(product_in[8]) );
  TBUF_X1 product_in_tri2_7_ ( .A(data_operandB[6]), .EN(n637), .Z(
        product_in[7]) );
  TBUF_X1 product_in_tri2_8_ ( .A(data_operandB[7]), .EN(n637), .Z(
        product_in[8]) );
  TBUF_X1 product_in_tri4_4_ ( .A(product_out[3]), .EN(n340), .Z(product_in[4]) );
  TBUF_X1 product_in_tri4_9_ ( .A(product_out[8]), .EN(n340), .Z(product_in[9]) );
  TBUF_X1 product_in_tri4_10_ ( .A(product_out[9]), .EN(n340), .Z(
        product_in[10]) );
  TBUF_X1 product_in_tri4_11_ ( .A(product_out[10]), .EN(n340), .Z(
        product_in[11]) );
  TBUF_X1 product_in_tri4_12_ ( .A(product_out[11]), .EN(n639), .Z(
        product_in[12]) );
  TBUF_X1 product_in_tri4_13_ ( .A(product_out[12]), .EN(n639), .Z(
        product_in[13]) );
  TBUF_X1 product_in_tri4_14_ ( .A(product_out[13]), .EN(n639), .Z(
        product_in[14]) );
  TBUF_X1 product_in_tri4_15_ ( .A(product_out[14]), .EN(n639), .Z(
        product_in[15]) );
  TBUF_X1 product_in_tri4_16_ ( .A(product_out[15]), .EN(n639), .Z(
        product_in[16]) );
  TBUF_X1 product_in_tri4_17_ ( .A(product_out[16]), .EN(n639), .Z(
        product_in[17]) );
  TBUF_X1 product_in_tri4_18_ ( .A(product_out[17]), .EN(n639), .Z(
        product_in[18]) );
  TBUF_X1 product_in_tri4_19_ ( .A(product_out[18]), .EN(n639), .Z(
        product_in[19]) );
  TBUF_X1 product_in_tri4_20_ ( .A(product_out[19]), .EN(n639), .Z(
        product_in[20]) );
  TBUF_X1 product_in_tri4_21_ ( .A(product_out[20]), .EN(n639), .Z(
        product_in[21]) );
  TBUF_X1 product_in_tri4_30_ ( .A(product_out[29]), .EN(n640), .Z(
        product_in[30]) );
  TBUF_X1 product_in_tri2_1_ ( .A(data_operandB[0]), .EN(n638), .Z(
        product_in[1]) );
  TBUF_X1 product_in_tri2_4_ ( .A(data_operandB[3]), .EN(n637), .Z(
        product_in[4]) );
  TBUF_X1 product_in_tri2_9_ ( .A(data_operandB[8]), .EN(n637), .Z(
        product_in[9]) );
  TBUF_X1 product_in_tri2_10_ ( .A(data_operandB[9]), .EN(n637), .Z(
        product_in[10]) );
  TBUF_X1 product_in_tri2_11_ ( .A(data_operandB[10]), .EN(n637), .Z(
        product_in[11]) );
  TBUF_X1 product_in_tri2_12_ ( .A(data_operandB[11]), .EN(n637), .Z(
        product_in[12]) );
  TBUF_X1 product_in_tri2_13_ ( .A(data_operandB[12]), .EN(n637), .Z(
        product_in[13]) );
  TBUF_X1 product_in_tri2_14_ ( .A(data_operandB[13]), .EN(n637), .Z(
        product_in[14]) );
  TBUF_X1 product_in_tri2_15_ ( .A(data_operandB[14]), .EN(n637), .Z(
        product_in[15]) );
  TBUF_X1 product_in_tri2_16_ ( .A(data_operandB[15]), .EN(n637), .Z(
        product_in[16]) );
  TBUF_X1 product_in_tri2_17_ ( .A(data_operandB[16]), .EN(n638), .Z(
        product_in[17]) );
  TBUF_X1 product_in_tri2_18_ ( .A(data_operandB[17]), .EN(n638), .Z(
        product_in[18]) );
  TBUF_X1 product_in_tri2_19_ ( .A(data_operandB[18]), .EN(n638), .Z(
        product_in[19]) );
  TBUF_X1 product_in_tri2_20_ ( .A(data_operandB[19]), .EN(n638), .Z(
        product_in[20]) );
  TBUF_X1 product_in_tri2_21_ ( .A(data_operandB[20]), .EN(n638), .Z(
        product_in[21]) );
  TBUF_X1 product_in_tri2_30_ ( .A(data_operandB[29]), .EN(n638), .Z(
        product_in[30]) );
  TBUF_X1 product_in_tri4_5_ ( .A(product_out[4]), .EN(n340), .Z(product_in[5]) );
  TBUF_X1 product_in_tri4_6_ ( .A(product_out[5]), .EN(n340), .Z(product_in[6]) );
  TBUF_X1 product_in_tri2_5_ ( .A(data_operandB[4]), .EN(n637), .Z(
        product_in[5]) );
  TBUF_X1 product_in_tri2_6_ ( .A(data_operandB[5]), .EN(n637), .Z(
        product_in[6]) );
  TBUF_X1 product_in_tri4_29_ ( .A(product_out[28]), .EN(n639), .Z(
        product_in[29]) );
  TBUF_X1 product_in_tri2_29_ ( .A(data_operandB[28]), .EN(n636), .Z(
        product_in[29]) );
  TBUF_X1 product_in_tri4_28_ ( .A(product_out[27]), .EN(n640), .Z(
        product_in[28]) );
  TBUF_X1 product_in_tri2_28_ ( .A(data_operandB[27]), .EN(n638), .Z(
        product_in[28]) );
  TBUF_X1 product_in_tri4_24_ ( .A(product_out[23]), .EN(n641), .Z(
        product_in[24]) );
  TBUF_X1 product_in_tri4_27_ ( .A(product_out[26]), .EN(n641), .Z(
        product_in[27]) );
  TBUF_X1 product_in_tri2_24_ ( .A(data_operandB[23]), .EN(n638), .Z(
        product_in[24]) );
  TBUF_X1 product_in_tri2_27_ ( .A(data_operandB[26]), .EN(n638), .Z(
        product_in[27]) );
  TBUF_X1 product_in_tri4_23_ ( .A(product_out[22]), .EN(n639), .Z(
        product_in[23]) );
  TBUF_X1 product_in_tri4_26_ ( .A(product_out[25]), .EN(n340), .Z(
        product_in[26]) );
  TBUF_X1 product_in_tri2_23_ ( .A(data_operandB[22]), .EN(n638), .Z(
        product_in[23]) );
  TBUF_X1 product_in_tri2_26_ ( .A(data_operandB[25]), .EN(n638), .Z(
        product_in[26]) );
  TBUF_X1 product_in_tri4_22_ ( .A(product_out[21]), .EN(n639), .Z(
        product_in[22]) );
  TBUF_X1 product_in_tri4_25_ ( .A(product_out[24]), .EN(n639), .Z(
        product_in[25]) );
  TBUF_X1 product_in_tri2_22_ ( .A(data_operandB[21]), .EN(n638), .Z(
        product_in[22]) );
  TBUF_X1 product_in_tri2_25_ ( .A(data_operandB[24]), .EN(n638), .Z(
        product_in[25]) );
  TBUF_X1 product_in_tri3_61_ ( .A(1'b0), .EN(n679), .Z(product_in[61]) );
  TBUF_X1 product_in_tri2_61_ ( .A(1'b0), .EN(n638), .Z(product_in[61]) );
  TBUF_X1 product_in_tri3_37_ ( .A(1'b0), .EN(n677), .Z(product_in[37]) );
  TBUF_X1 product_in_tri3_39_ ( .A(1'b0), .EN(n677), .Z(product_in[39]) );
  TBUF_X1 product_in_tri3_40_ ( .A(1'b0), .EN(n677), .Z(product_in[40]) );
  TBUF_X1 product_in_tri3_42_ ( .A(1'b0), .EN(n677), .Z(product_in[42]) );
  TBUF_X1 product_in_tri3_45_ ( .A(1'b0), .EN(n677), .Z(product_in[45]) );
  TBUF_X1 product_in_tri3_47_ ( .A(1'b0), .EN(n677), .Z(product_in[47]) );
  TBUF_X1 product_in_tri3_48_ ( .A(1'b0), .EN(n677), .Z(product_in[48]) );
  TBUF_X1 product_in_tri3_50_ ( .A(1'b0), .EN(n679), .Z(product_in[50]) );
  TBUF_X1 product_in_tri3_53_ ( .A(1'b0), .EN(n679), .Z(product_in[53]) );
  TBUF_X1 product_in_tri3_55_ ( .A(1'b0), .EN(n679), .Z(product_in[55]) );
  TBUF_X1 product_in_tri3_56_ ( .A(1'b0), .EN(n679), .Z(product_in[56]) );
  TBUF_X1 product_in_tri3_58_ ( .A(1'b0), .EN(n679), .Z(product_in[58]) );
  TBUF_X1 product_in_tri2_37_ ( .A(1'b0), .EN(n635), .Z(product_in[37]) );
  TBUF_X1 product_in_tri2_39_ ( .A(1'b0), .EN(n635), .Z(product_in[39]) );
  TBUF_X1 product_in_tri2_40_ ( .A(1'b0), .EN(n635), .Z(product_in[40]) );
  TBUF_X1 product_in_tri2_42_ ( .A(1'b0), .EN(n635), .Z(product_in[42]) );
  TBUF_X1 product_in_tri2_45_ ( .A(1'b0), .EN(n636), .Z(product_in[45]) );
  TBUF_X1 product_in_tri2_47_ ( .A(1'b0), .EN(n636), .Z(product_in[47]) );
  TBUF_X1 product_in_tri2_48_ ( .A(1'b0), .EN(n636), .Z(product_in[48]) );
  TBUF_X1 product_in_tri2_50_ ( .A(1'b0), .EN(n636), .Z(product_in[50]) );
  TBUF_X1 product_in_tri2_53_ ( .A(1'b0), .EN(n636), .Z(product_in[53]) );
  TBUF_X1 product_in_tri2_55_ ( .A(1'b0), .EN(n636), .Z(product_in[55]) );
  TBUF_X1 product_in_tri2_56_ ( .A(1'b0), .EN(n637), .Z(product_in[56]) );
  TBUF_X1 product_in_tri2_58_ ( .A(1'b0), .EN(n636), .Z(product_in[58]) );
  TBUF_X1 product_in_tri3_35_ ( .A(1'b0), .EN(n678), .Z(product_in[35]) );
  TBUF_X1 product_in_tri3_60_ ( .A(1'b0), .EN(n679), .Z(product_in[60]) );
  TBUF_X1 product_in_tri2_35_ ( .A(1'b0), .EN(n635), .Z(product_in[35]) );
  TBUF_X1 product_in_tri2_60_ ( .A(1'b0), .EN(n637), .Z(product_in[60]) );
  TBUF_X1 product_in_tri3_36_ ( .A(1'b0), .EN(n677), .Z(product_in[36]) );
  TBUF_X1 product_in_tri3_38_ ( .A(1'b0), .EN(n678), .Z(product_in[38]) );
  TBUF_X1 product_in_tri3_41_ ( .A(1'b0), .EN(n678), .Z(product_in[41]) );
  TBUF_X1 product_in_tri3_43_ ( .A(1'b0), .EN(n678), .Z(product_in[43]) );
  TBUF_X1 product_in_tri3_44_ ( .A(1'b0), .EN(n679), .Z(product_in[44]) );
  TBUF_X1 product_in_tri3_46_ ( .A(1'b0), .EN(n679), .Z(product_in[46]) );
  TBUF_X1 product_in_tri3_49_ ( .A(1'b0), .EN(n679), .Z(product_in[49]) );
  TBUF_X1 product_in_tri3_51_ ( .A(1'b0), .EN(n679), .Z(product_in[51]) );
  TBUF_X1 product_in_tri3_52_ ( .A(1'b0), .EN(n679), .Z(product_in[52]) );
  TBUF_X1 product_in_tri3_54_ ( .A(1'b0), .EN(n679), .Z(product_in[54]) );
  TBUF_X1 product_in_tri3_57_ ( .A(1'b0), .EN(n679), .Z(product_in[57]) );
  TBUF_X1 product_in_tri3_59_ ( .A(1'b0), .EN(n679), .Z(product_in[59]) );
  TBUF_X1 product_in_tri2_36_ ( .A(1'b0), .EN(n635), .Z(product_in[36]) );
  TBUF_X1 product_in_tri2_38_ ( .A(1'b0), .EN(n635), .Z(product_in[38]) );
  TBUF_X1 product_in_tri2_41_ ( .A(1'b0), .EN(n635), .Z(product_in[41]) );
  TBUF_X1 product_in_tri2_43_ ( .A(1'b0), .EN(n635), .Z(product_in[43]) );
  TBUF_X1 product_in_tri2_44_ ( .A(1'b0), .EN(n636), .Z(product_in[44]) );
  TBUF_X1 product_in_tri2_46_ ( .A(1'b0), .EN(n636), .Z(product_in[46]) );
  TBUF_X1 product_in_tri2_49_ ( .A(1'b0), .EN(n636), .Z(product_in[49]) );
  TBUF_X1 product_in_tri2_51_ ( .A(1'b0), .EN(n636), .Z(product_in[51]) );
  TBUF_X1 product_in_tri2_52_ ( .A(1'b0), .EN(n636), .Z(product_in[52]) );
  TBUF_X1 product_in_tri2_54_ ( .A(1'b0), .EN(n636), .Z(product_in[54]) );
  TBUF_X1 product_in_tri2_57_ ( .A(1'b0), .EN(n638), .Z(product_in[57]) );
  TBUF_X1 product_in_tri2_59_ ( .A(1'b0), .EN(n637), .Z(product_in[59]) );
  TBUF_X1 product_in_tri2_64_ ( .A(1'b0), .EN(n635), .Z(product_in[64]) );
  TBUF_X1 product_in_tri3_33_ ( .A(1'b0), .EN(n679), .Z(product_in[33]) );
  TBUF_X1 product_in_tri2_33_ ( .A(1'b0), .EN(n635), .Z(product_in[33]) );
  TBUF_X1 product_in_tri4_0_ ( .A(1'b0), .EN(n340), .Z(product_in[0]) );
  TBUF_X1 product_in_tri3_0_ ( .A(1'b0), .EN(n677), .Z(product_in[0]) );
  TBUF_X1 product_in_tri2_0_ ( .A(1'b0), .EN(n636), .Z(product_in[0]) );
  TBUF_X1 product_in_tri2_3_ ( .A(data_operandB[2]), .EN(n638), .Z(
        product_in[3]) );
  TBUF_X1 product_in_tri2_2_ ( .A(data_operandB[1]), .EN(n461), .Z(
        product_in[2]) );
  TBUF_X1 product_in_tri4_31_ ( .A(product_out[30]), .EN(n641), .Z(
        product_in[31]) );
  TBUF_X1 product_in_tri2_31_ ( .A(data_operandB[30]), .EN(n637), .Z(
        product_in[31]) );
  TBUF_X1 product_in_tri4_32_ ( .A(product_out[31]), .EN(n639), .Z(
        product_in[32]) );
  TBUF_X1 product_in_tri3_34_ ( .A(1'b0), .EN(n677), .Z(product_in[34]) );
  TBUF_X1 product_in_tri2_34_ ( .A(1'b0), .EN(n635), .Z(product_in[34]) );
  TBUF_X1 product_in_tri2_32_ ( .A(data_operandB[31]), .EN(n636), .Z(
        product_in[32]) );
  TBUF_X1 product_in_tri3_7_ ( .A(n213), .EN(n679), .Z(product_in[7]) );
  TBUF_X1 product_in_tri3_8_ ( .A(n212), .EN(n678), .Z(product_in[8]) );
  TBUF_X1 product_in_tri_7_ ( .A(product_out[9]), .EN(n654), .Z(product_in[7])
         );
  TBUF_X1 product_in_tri_8_ ( .A(product_out[10]), .EN(n654), .Z(product_in[8]) );
  TBUF_X1 product_in_tri3_1_ ( .A(n367), .EN(n679), .Z(product_in[1]) );
  TBUF_X1 product_in_tri3_4_ ( .A(n370), .EN(n679), .Z(product_in[4]) );
  TBUF_X1 product_in_tri_1_ ( .A(product_out[3]), .EN(n654), .Z(product_in[1])
         );
  TBUF_X1 product_in_tri_4_ ( .A(product_out[6]), .EN(n654), .Z(product_in[4])
         );
  TBUF_X1 product_in_tri_9_ ( .A(product_out[11]), .EN(n654), .Z(product_in[9]) );
  TBUF_X1 product_in_tri_10_ ( .A(product_out[12]), .EN(n654), .Z(
        product_in[10]) );
  TBUF_X1 product_in_tri_11_ ( .A(product_out[13]), .EN(n654), .Z(
        product_in[11]) );
  TBUF_X1 product_in_tri_12_ ( .A(product_out[14]), .EN(n653), .Z(
        product_in[12]) );
  TBUF_X1 product_in_tri_13_ ( .A(product_out[15]), .EN(n653), .Z(
        product_in[13]) );
  TBUF_X1 product_in_tri_14_ ( .A(product_out[16]), .EN(n653), .Z(
        product_in[14]) );
  TBUF_X1 product_in_tri_15_ ( .A(product_out[17]), .EN(n653), .Z(
        product_in[15]) );
  TBUF_X1 product_in_tri_16_ ( .A(product_out[18]), .EN(n653), .Z(
        product_in[16]) );
  TBUF_X1 product_in_tri_17_ ( .A(product_out[19]), .EN(n653), .Z(
        product_in[17]) );
  TBUF_X1 product_in_tri_18_ ( .A(product_out[20]), .EN(n653), .Z(
        product_in[18]) );
  TBUF_X1 product_in_tri_19_ ( .A(product_out[21]), .EN(n653), .Z(
        product_in[19]) );
  TBUF_X1 product_in_tri_20_ ( .A(product_out[22]), .EN(n653), .Z(
        product_in[20]) );
  TBUF_X1 product_in_tri_21_ ( .A(product_out[23]), .EN(n653), .Z(
        product_in[21]) );
  TBUF_X1 product_in_tri_30_ ( .A(product_out[32]), .EN(n630), .Z(
        product_in[30]) );
  TBUF_X1 product_in_tri3_13_ ( .A(n379), .EN(n678), .Z(product_in[13]) );
  TBUF_X1 product_in_tri3_14_ ( .A(n380), .EN(n679), .Z(product_in[14]) );
  TBUF_X1 product_in_tri3_15_ ( .A(n381), .EN(n678), .Z(product_in[15]) );
  TBUF_X1 product_in_tri3_16_ ( .A(n382), .EN(n678), .Z(product_in[16]) );
  TBUF_X1 product_in_tri3_9_ ( .A(n210), .EN(n679), .Z(product_in[9]) );
  TBUF_X1 product_in_tri3_10_ ( .A(n209), .EN(n678), .Z(product_in[10]) );
  TBUF_X1 product_in_tri3_11_ ( .A(n377), .EN(n679), .Z(product_in[11]) );
  TBUF_X1 product_in_tri3_12_ ( .A(n378), .EN(n678), .Z(product_in[12]) );
  TBUF_X1 product_in_tri3_17_ ( .A(n383), .EN(n678), .Z(product_in[17]) );
  TBUF_X1 product_in_tri3_18_ ( .A(n384), .EN(n678), .Z(product_in[18]) );
  TBUF_X1 product_in_tri3_19_ ( .A(n385), .EN(n678), .Z(product_in[19]) );
  TBUF_X1 product_in_tri3_20_ ( .A(n386), .EN(n678), .Z(product_in[20]) );
  TBUF_X1 product_in_tri3_21_ ( .A(n198), .EN(n678), .Z(product_in[21]) );
  TBUF_X1 product_in_tri3_5_ ( .A(n371), .EN(n679), .Z(product_in[5]) );
  TBUF_X1 product_in_tri3_6_ ( .A(n214), .EN(n678), .Z(product_in[6]) );
  TBUF_X1 product_in_tri_5_ ( .A(product_out[7]), .EN(n654), .Z(product_in[5])
         );
  TBUF_X1 product_in_tri_6_ ( .A(product_out[8]), .EN(n654), .Z(product_in[6])
         );
  TBUF_X1 product_in_tri_29_ ( .A(product_out[31]), .EN(n618), .Z(
        product_in[29]) );
  TBUF_X1 product_in_tri_28_ ( .A(product_out[30]), .EN(n630), .Z(
        product_in[28]) );
  TBUF_X1 product_in_tri_24_ ( .A(product_out[26]), .EN(n653), .Z(
        product_in[24]) );
  TBUF_X1 product_in_tri_27_ ( .A(product_out[29]), .EN(n618), .Z(
        product_in[27]) );
  TBUF_X1 product_in_tri_23_ ( .A(product_out[25]), .EN(n653), .Z(
        product_in[23]) );
  TBUF_X1 product_in_tri_26_ ( .A(product_out[28]), .EN(n630), .Z(
        product_in[26]) );
  TBUF_X1 product_in_tri3_23_ ( .A(n196), .EN(n678), .Z(product_in[23]) );
  TBUF_X1 product_in_tri_22_ ( .A(product_out[24]), .EN(n653), .Z(
        product_in[22]) );
  TBUF_X1 product_in_tri_25_ ( .A(product_out[27]), .EN(n618), .Z(
        product_in[25]) );
  TBUF_X1 product_in_tri3_22_ ( .A(n197), .EN(n678), .Z(product_in[22]) );
  TBUF_X1 product_in_tri4_37_ ( .A(adder_out[4]), .EN(n640), .Z(product_in[37]) );
  TBUF_X1 product_in_tri_39_ ( .A(adder_out[8]), .EN(n656), .Z(product_in[39])
         );
  TBUF_X1 product_in_tri_40_ ( .A(adder_out[9]), .EN(n656), .Z(product_in[40])
         );
  TBUF_X1 product_in_tri4_42_ ( .A(adder_out[9]), .EN(n640), .Z(product_in[42]) );
  TBUF_X1 product_in_tri4_39_ ( .A(adder_out[6]), .EN(n640), .Z(product_in[39]) );
  TBUF_X1 product_in_tri4_40_ ( .A(adder_out[7]), .EN(n640), .Z(product_in[40]) );
  TBUF_X1 product_in_tri_37_ ( .A(adder_out[6]), .EN(n656), .Z(product_in[37])
         );
  TBUF_X1 product_in_tri_42_ ( .A(adder_out[11]), .EN(n656), .Z(product_in[42]) );
  TBUF_X1 product_in_tri4_45_ ( .A(adder_out[12]), .EN(n640), .Z(
        product_in[45]) );
  TBUF_X1 product_in_tri4_47_ ( .A(adder_out[14]), .EN(n640), .Z(
        product_in[47]) );
  TBUF_X1 product_in_tri_45_ ( .A(adder_out[14]), .EN(n656), .Z(product_in[45]) );
  TBUF_X1 product_in_tri4_48_ ( .A(adder_out[15]), .EN(n641), .Z(
        product_in[48]) );
  TBUF_X1 product_in_tri_47_ ( .A(adder_out[16]), .EN(n656), .Z(product_in[47]) );
  TBUF_X1 product_in_tri4_50_ ( .A(adder_out[17]), .EN(n641), .Z(
        product_in[50]) );
  TBUF_X1 product_in_tri_48_ ( .A(adder_out[17]), .EN(n655), .Z(product_in[48]) );
  TBUF_X1 product_in_tri_50_ ( .A(adder_out[19]), .EN(n655), .Z(product_in[50]) );
  TBUF_X1 product_in_tri4_53_ ( .A(adder_out[20]), .EN(n641), .Z(
        product_in[53]) );
  TBUF_X1 product_in_tri4_35_ ( .A(adder_out[2]), .EN(n340), .Z(product_in[35]) );
  TBUF_X1 product_in_tri_35_ ( .A(adder_out[4]), .EN(n656), .Z(product_in[35])
         );
  TBUF_X1 product_in_tri4_36_ ( .A(adder_out[3]), .EN(n640), .Z(product_in[36]) );
  TBUF_X1 product_in_tri4_41_ ( .A(adder_out[8]), .EN(n640), .Z(product_in[41]) );
  TBUF_X1 product_in_tri4_43_ ( .A(adder_out[10]), .EN(n640), .Z(
        product_in[43]) );
  TBUF_X1 product_in_tri_41_ ( .A(adder_out[10]), .EN(n656), .Z(product_in[41]) );
  TBUF_X1 product_in_tri4_38_ ( .A(adder_out[5]), .EN(n640), .Z(product_in[38]) );
  TBUF_X1 product_in_tri_36_ ( .A(adder_out[5]), .EN(n656), .Z(product_in[36])
         );
  TBUF_X1 product_in_tri_38_ ( .A(adder_out[7]), .EN(n656), .Z(product_in[38])
         );
  TBUF_X1 product_in_tri4_44_ ( .A(adder_out[11]), .EN(n640), .Z(
        product_in[44]) );
  TBUF_X1 product_in_tri_43_ ( .A(adder_out[12]), .EN(n656), .Z(product_in[43]) );
  TBUF_X1 product_in_tri4_46_ ( .A(adder_out[13]), .EN(n640), .Z(
        product_in[46]) );
  TBUF_X1 product_in_tri_44_ ( .A(adder_out[13]), .EN(n656), .Z(product_in[44]) );
  TBUF_X1 product_in_tri_46_ ( .A(adder_out[15]), .EN(n656), .Z(product_in[46]) );
  TBUF_X1 product_in_tri4_49_ ( .A(adder_out[16]), .EN(n641), .Z(
        product_in[49]) );
  TBUF_X1 product_in_tri4_51_ ( .A(adder_out[18]), .EN(n641), .Z(
        product_in[51]) );
  TBUF_X1 product_in_tri_49_ ( .A(adder_out[18]), .EN(n655), .Z(product_in[49]) );
  TBUF_X1 product_in_tri4_52_ ( .A(adder_out[19]), .EN(n641), .Z(
        product_in[52]) );
  TBUF_X1 product_in_tri_51_ ( .A(adder_out[20]), .EN(n655), .Z(product_in[51]) );
  TBUF_X1 product_in_tri3_3_ ( .A(n369), .EN(n679), .Z(product_in[3]) );
  TBUF_X1 product_in_tri_3_ ( .A(product_out[5]), .EN(n654), .Z(product_in[3])
         );
  TBUF_X1 product_in_tri3_2_ ( .A(n368), .EN(n678), .Z(product_in[2]) );
  TBUF_X1 product_in_tri_2_ ( .A(product_out[4]), .EN(n654), .Z(product_in[2])
         );
  TBUF_X1 product_in_tri4_34_ ( .A(adder_out[1]), .EN(n340), .Z(product_in[34]) );
  TBUF_X1 product_in_tri3_30_ ( .A(n396), .EN(n677), .Z(product_in[30]) );
  TBUF_X1 product_in_tri4_1_ ( .A(n366), .EN(n340), .Z(product_in[1]) );
  TBUF_X1 product_in_tri3_29_ ( .A(n395), .EN(n678), .Z(product_in[29]) );
  TBUF_X1 product_in_tri3_28_ ( .A(n394), .EN(n678), .Z(product_in[28]) );
  TBUF_X1 product_in_tri3_24_ ( .A(n390), .EN(n678), .Z(product_in[24]) );
  TBUF_X1 product_in_tri3_27_ ( .A(n393), .EN(n678), .Z(product_in[27]) );
  TBUF_X1 product_in_tri3_26_ ( .A(n392), .EN(n678), .Z(product_in[26]) );
  TBUF_X1 product_in_tri3_25_ ( .A(n391), .EN(n678), .Z(product_in[25]) );
  TBUF_X1 product_in_tri4_61_ ( .A(adder_out[28]), .EN(n340), .Z(
        product_in[61]) );
  TBUF_X1 product_in_tri_61_ ( .A(adder_out[30]), .EN(n654), .Z(product_in[61]) );
  TBUF_X1 product_in_tri4_55_ ( .A(adder_out[22]), .EN(n641), .Z(
        product_in[55]) );
  TBUF_X1 product_in_tri_53_ ( .A(adder_out[22]), .EN(n655), .Z(product_in[53]) );
  TBUF_X1 product_in_tri4_56_ ( .A(adder_out[23]), .EN(n641), .Z(
        product_in[56]) );
  TBUF_X1 product_in_tri_55_ ( .A(adder_out[24]), .EN(n655), .Z(product_in[55]) );
  TBUF_X1 product_in_tri4_58_ ( .A(adder_out[25]), .EN(n641), .Z(
        product_in[58]) );
  TBUF_X1 product_in_tri_56_ ( .A(adder_out[25]), .EN(n655), .Z(product_in[56]) );
  TBUF_X1 product_in_tri_58_ ( .A(adder_out[27]), .EN(n655), .Z(product_in[58]) );
  TBUF_X1 product_in_tri4_60_ ( .A(adder_out[27]), .EN(n340), .Z(
        product_in[60]) );
  TBUF_X1 product_in_tri_60_ ( .A(n613), .EN(n655), .Z(product_in[60]) );
  TBUF_X1 product_in_tri4_54_ ( .A(adder_out[21]), .EN(n641), .Z(
        product_in[54]) );
  TBUF_X1 product_in_tri_52_ ( .A(adder_out[21]), .EN(n655), .Z(product_in[52]) );
  TBUF_X1 product_in_tri_54_ ( .A(adder_out[23]), .EN(n655), .Z(product_in[54]) );
  TBUF_X1 product_in_tri4_57_ ( .A(adder_out[24]), .EN(n641), .Z(
        product_in[57]) );
  TBUF_X1 product_in_tri4_59_ ( .A(adder_out[26]), .EN(n641), .Z(
        product_in[59]) );
  TBUF_X1 product_in_tri_57_ ( .A(adder_out[26]), .EN(n655), .Z(product_in[57]) );
  TBUF_X1 product_in_tri_59_ ( .A(adder_out[28]), .EN(n655), .Z(product_in[59]) );
  TBUF_X1 product_in_tri3_31_ ( .A(n397), .EN(n677), .Z(product_in[31]) );
  TBUF_X1 product_in_tri3_32_ ( .A(n187), .EN(n677), .Z(product_in[32]) );
  INV_X1 U712 ( .A(n643), .ZN(n650) );
  BUF_X1 U713 ( .A(n643), .Z(n660) );
  BUF_X1 U714 ( .A(n644), .Z(n664) );
  BUF_X1 U715 ( .A(n644), .Z(n662) );
  BUF_X1 U716 ( .A(op_mult), .Z(n647) );
  CLKBUF_X1 U717 ( .A(n643), .Z(n661) );
  BUF_X1 U718 ( .A(op_mult), .Z(n621) );
  BUF_X2 U719 ( .A(ctrl_DIV), .Z(n673) );
  OR2_X1 U720 ( .A1(n339), .A2(n522), .ZN(n611) );
  CLKBUF_X1 U721 ( .A(operandA[0]), .Z(n627) );
  CLKBUF_X1 U722 ( .A(op_mult), .Z(n645) );
  BUF_X1 U723 ( .A(n363), .Z(n626) );
  CLKBUF_X1 U724 ( .A(operandA[4]), .Z(n612) );
  CLKBUF_X1 U725 ( .A(product_in[63]), .Z(n631) );
  BUF_X1 U726 ( .A(op_mult), .Z(n646) );
  BUF_X1 U727 ( .A(adder_out[29]), .Z(n613) );
  BUF_X1 U728 ( .A(ctrl_DIV), .Z(n614) );
  BUF_X1 U729 ( .A(ctrl_MULT), .Z(n615) );
  MUX2_X1 U730 ( .A(product_out[2]), .B(data_operandA[1]), .S(ctrl_DIV), .Z(
        n616) );
  INV_X1 U731 ( .A(n616), .ZN(n580) );
  MUX2_X1 U732 ( .A(data_operandA[30]), .B(sign_fixed[30]), .S(
        data_operandA[31]), .Z(n397) );
  MUX2_X1 U733 ( .A(product_out[1]), .B(data_operandA[0]), .S(ctrl_DIV), .Z(
        n617) );
  INV_X1 U734 ( .A(n617), .ZN(n579) );
  INV_X1 U735 ( .A(n665), .ZN(n618) );
  BUF_X1 U736 ( .A(n645), .Z(n665) );
  CLKBUF_X1 U737 ( .A(product_out[1]), .Z(n619) );
  AND2_X1 U738 ( .A1(data_operandA[31]), .A2(sign_fixed[31]), .ZN(n187) );
  CLKBUF_X1 U739 ( .A(operandA[2]), .Z(n620) );
  INV_X1 U740 ( .A(n567), .ZN(n622) );
  CLKBUF_X1 U741 ( .A(adder_out[31]), .Z(n623) );
  CLKBUF_X1 U742 ( .A(product_out[2]), .Z(n624) );
  CLKBUF_X3 U743 ( .A(n621), .Z(n668) );
  CLKBUF_X1 U744 ( .A(operandA_shift_0_), .Z(n629) );
  AND2_X1 U745 ( .A1(product_in[62]), .A2(n660), .ZN(n625) );
  CLKBUF_X1 U746 ( .A(product_in[62]), .Z(n628) );
  INV_X2 U747 ( .A(n644), .ZN(n651) );
  CLKBUF_X1 U748 ( .A(n642), .Z(n657) );
  CLKBUF_X1 U749 ( .A(n642), .Z(n658) );
  CLKBUF_X1 U750 ( .A(n647), .Z(n666) );
  INV_X2 U751 ( .A(n646), .ZN(n649) );
  INV_X2 U752 ( .A(n671), .ZN(n676) );
  BUF_X1 U753 ( .A(ctrl_DIV), .Z(n674) );
  INV_X1 U754 ( .A(n668), .ZN(n656) );
  CLKBUF_X1 U755 ( .A(n649), .Z(n630) );
  CLKBUF_X1 U756 ( .A(n644), .Z(n663) );
  BUF_X1 U757 ( .A(n642), .Z(n659) );
  CLKBUF_X1 U758 ( .A(n647), .Z(n667) );
  INV_X1 U759 ( .A(n611), .ZN(n633) );
  INV_X1 U760 ( .A(n611), .ZN(n632) );
  CLKBUF_X1 U761 ( .A(n645), .Z(n642) );
  BUF_X1 U762 ( .A(n611), .Z(n634) );
  INV_X1 U763 ( .A(data_operandA[31]), .ZN(n680) );
  INV_X1 U764 ( .A(data_operandA[31]), .ZN(n681) );
  INV_X1 U765 ( .A(data_resultRDY), .ZN(n365) );
  INV_X1 U766 ( .A(n674), .ZN(n675) );
  OAI22_X1 U767 ( .A1(n649), .A2(n413), .B1(n658), .B2(n412), .ZN(n_2_net__5_)
         );
  OAI22_X1 U768 ( .A1(n630), .A2(n412), .B1(n658), .B2(n411), .ZN(n_2_net__4_)
         );
  OAI22_X1 U769 ( .A1(n649), .A2(n415), .B1(n657), .B2(n414), .ZN(n_2_net__7_)
         );
  OAI22_X1 U770 ( .A1(n651), .A2(n414), .B1(n657), .B2(n413), .ZN(n_2_net__6_)
         );
  OAI22_X1 U771 ( .A1(n649), .A2(n411), .B1(n658), .B2(n410), .ZN(n_2_net__3_)
         );
  OAI22_X1 U772 ( .A1(n650), .A2(n410), .B1(n659), .B2(n409), .ZN(n_2_net__2_)
         );
  OAI22_X1 U773 ( .A1(n651), .A2(n408), .B1(n663), .B2(n407), .ZN(n_2_net__0_)
         );
  OAI22_X1 U774 ( .A1(n650), .A2(n409), .B1(n667), .B2(n408), .ZN(n_2_net__1_)
         );
  OAI22_X1 U775 ( .A1(n665), .A2(n458), .B1(n648), .B2(n448), .ZN(n_1_net__5_)
         );
  OAI22_X1 U776 ( .A1(n665), .A2(n457), .B1(n648), .B2(n447), .ZN(n_1_net__6_)
         );
  OAI22_X1 U777 ( .A1(n665), .A2(n454), .B1(n648), .B2(n444), .ZN(n_1_net__9_)
         );
  INV_X1 U778 ( .A(n556), .ZN(n341) );
  OAI22_X1 U779 ( .A1(n666), .A2(n456), .B1(n648), .B2(n446), .ZN(n_1_net__7_)
         );
  INV_X1 U780 ( .A(n577), .ZN(n362) );
  INV_X1 U781 ( .A(n573), .ZN(n358) );
  INV_X1 U782 ( .A(n574), .ZN(n359) );
  INV_X1 U783 ( .A(n575), .ZN(n360) );
  INV_X1 U784 ( .A(n559), .ZN(n344) );
  OAI22_X1 U785 ( .A1(n665), .A2(n455), .B1(n648), .B2(n445), .ZN(n_1_net__8_)
         );
  INV_X1 U786 ( .A(n572), .ZN(n357) );
  INV_X1 U787 ( .A(n576), .ZN(n361) );
  INV_X1 U788 ( .A(n673), .ZN(n677) );
  OAI22_X1 U789 ( .A1(n650), .A2(n416), .B1(n657), .B2(n415), .ZN(n_2_net__8_)
         );
  OAI22_X1 U790 ( .A1(n651), .A2(n424), .B1(n662), .B2(n423), .ZN(n_2_net__16_) );
  OAI22_X1 U791 ( .A1(n651), .A2(n421), .B1(n663), .B2(n420), .ZN(n_2_net__13_) );
  OAI22_X1 U792 ( .A1(n618), .A2(n420), .B1(n662), .B2(n419), .ZN(n_2_net__12_) );
  OAI22_X1 U793 ( .A1(n650), .A2(n418), .B1(n663), .B2(n417), .ZN(n_2_net__10_) );
  OAI22_X1 U794 ( .A1(n651), .A2(n428), .B1(n661), .B2(n427), .ZN(n_2_net__20_) );
  OAI22_X1 U795 ( .A1(n650), .A2(n426), .B1(n664), .B2(n425), .ZN(n_2_net__18_) );
  OAI22_X1 U796 ( .A1(n651), .A2(n429), .B1(n661), .B2(n428), .ZN(n_2_net__21_) );
  OAI22_X1 U797 ( .A1(n648), .A2(n437), .B1(n659), .B2(n436), .ZN(n_2_net__29_) );
  OAI22_X1 U798 ( .A1(n651), .A2(n436), .B1(n659), .B2(n435), .ZN(n_2_net__28_) );
  OAI22_X1 U799 ( .A1(n618), .A2(n434), .B1(n660), .B2(n433), .ZN(n_2_net__26_) );
  OAI22_X1 U800 ( .A1(n651), .A2(n432), .B1(n660), .B2(n431), .ZN(n_2_net__24_) );
  OAI22_X1 U801 ( .A1(n650), .A2(n431), .B1(n661), .B2(n430), .ZN(n_2_net__23_) );
  OAI22_X1 U802 ( .A1(n651), .A2(n423), .B1(n662), .B2(n422), .ZN(n_2_net__15_) );
  OAI22_X1 U803 ( .A1(n650), .A2(n439), .B1(n658), .B2(n438), .ZN(n_2_net__31_) );
  OAI22_X1 U804 ( .A1(n650), .A2(n417), .B1(n657), .B2(n416), .ZN(n_2_net__9_)
         );
  OAI22_X1 U805 ( .A1(n630), .A2(n425), .B1(n662), .B2(n424), .ZN(n_2_net__17_) );
  OAI22_X1 U806 ( .A1(n651), .A2(n430), .B1(n661), .B2(n429), .ZN(n_2_net__22_) );
  OAI22_X1 U807 ( .A1(n650), .A2(n422), .B1(n663), .B2(n421), .ZN(n_2_net__14_) );
  OAI22_X1 U808 ( .A1(n651), .A2(n419), .B1(n660), .B2(n418), .ZN(n_2_net__11_) );
  OAI22_X1 U809 ( .A1(n651), .A2(n427), .B1(n664), .B2(n426), .ZN(n_2_net__19_) );
  OAI22_X1 U810 ( .A1(n650), .A2(n435), .B1(n660), .B2(n434), .ZN(n_2_net__27_) );
  OAI22_X1 U811 ( .A1(n650), .A2(n438), .B1(n659), .B2(n437), .ZN(n_2_net__30_) );
  OAI22_X1 U812 ( .A1(n650), .A2(n433), .B1(n660), .B2(n432), .ZN(n_2_net__25_) );
  OAI22_X1 U813 ( .A1(n680), .A2(n389), .B1(data_operandA[31]), .B2(n441), 
        .ZN(n196) );
  OAI22_X1 U814 ( .A1(n680), .A2(n388), .B1(data_operandA[31]), .B2(n442), 
        .ZN(n197) );
  OAI22_X1 U815 ( .A1(n680), .A2(n387), .B1(data_operandA[31]), .B2(n443), 
        .ZN(n198) );
  OAI22_X1 U816 ( .A1(n680), .A2(n376), .B1(data_operandA[31]), .B2(n444), 
        .ZN(n209) );
  OAI22_X1 U817 ( .A1(n680), .A2(n375), .B1(data_operandA[31]), .B2(n445), 
        .ZN(n210) );
  OAI22_X1 U818 ( .A1(n680), .A2(n374), .B1(data_operandA[31]), .B2(n446), 
        .ZN(n212) );
  OAI22_X1 U819 ( .A1(n680), .A2(n373), .B1(data_operandA[31]), .B2(n447), 
        .ZN(n213) );
  OAI22_X1 U820 ( .A1(n680), .A2(n372), .B1(data_operandA[31]), .B2(n448), 
        .ZN(n214) );
  OAI22_X1 U821 ( .A1(n664), .A2(n453), .B1(n648), .B2(n443), .ZN(n_1_net__20_) );
  OAI22_X1 U822 ( .A1(n664), .A2(n452), .B1(n618), .B2(n442), .ZN(n_1_net__21_) );
  INV_X1 U823 ( .A(n571), .ZN(n356) );
  INV_X1 U824 ( .A(n568), .ZN(n353) );
  INV_X1 U825 ( .A(n569), .ZN(n354) );
  INV_X1 U826 ( .A(n560), .ZN(n345) );
  INV_X1 U827 ( .A(n558), .ZN(n343) );
  INV_X1 U828 ( .A(n564), .ZN(n349) );
  INV_X1 U829 ( .A(n562), .ZN(n347) );
  INV_X1 U830 ( .A(sign_fixed[22]), .ZN(n389) );
  INV_X1 U831 ( .A(sign_fixed[9]), .ZN(n376) );
  INV_X1 U832 ( .A(sign_fixed[6]), .ZN(n373) );
  OAI22_X1 U833 ( .A1(n664), .A2(n451), .B1(n648), .B2(n441), .ZN(n_1_net__22_) );
  OAI22_X1 U834 ( .A1(n664), .A2(n449), .B1(n648), .B2(n680), .ZN(n_1_net__31_) );
  INV_X1 U835 ( .A(n566), .ZN(n351) );
  INV_X1 U836 ( .A(n565), .ZN(n350) );
  INV_X1 U837 ( .A(n563), .ZN(n348) );
  INV_X1 U838 ( .A(n561), .ZN(n346) );
  INV_X1 U839 ( .A(n570), .ZN(n355) );
  INV_X1 U840 ( .A(n674), .ZN(n678) );
  INV_X1 U841 ( .A(n674), .ZN(n679) );
  BUF_X1 U842 ( .A(n461), .Z(n638) );
  BUF_X1 U843 ( .A(n461), .Z(n637) );
  BUF_X1 U844 ( .A(n461), .Z(n636) );
  BUF_X1 U845 ( .A(n461), .Z(n635) );
  BUF_X1 U846 ( .A(n340), .Z(n641) );
  BUF_X1 U847 ( .A(n340), .Z(n640) );
  BUF_X1 U848 ( .A(n340), .Z(n639) );
  NOR4_X1 U849 ( .A1(n540), .A2(n541), .A3(n542), .A4(n543), .ZN(n539) );
  NAND4_X1 U850 ( .A1(n415), .A2(n416), .A3(n417), .A4(n418), .ZN(n541) );
  NAND4_X1 U851 ( .A1(n419), .A2(n420), .A3(n421), .A4(n422), .ZN(n540) );
  NAND4_X1 U852 ( .A1(n407), .A2(n408), .A3(n409), .A4(n410), .ZN(n543) );
  OAI22_X1 U853 ( .A1(n398), .A2(n611), .B1(n633), .B2(n407), .ZN(
        data_result[31]) );
  AOI211_X1 U854 ( .C1(n526), .C2(n527), .A(n522), .B(data_result[31]), .ZN(
        n525) );
  NOR4_X1 U855 ( .A1(n532), .A2(n533), .A3(n534), .A4(n535), .ZN(n526) );
  NOR4_X1 U856 ( .A1(n528), .A2(n529), .A3(n530), .A4(n531), .ZN(n527) );
  OAI22_X1 U857 ( .A1(n372), .A2(n634), .B1(n632), .B2(n399), .ZN(
        data_result[5]) );
  OAI22_X1 U858 ( .A1(n373), .A2(n634), .B1(n633), .B2(n400), .ZN(
        data_result[6]) );
  OAI22_X1 U859 ( .A1(n374), .A2(n611), .B1(n632), .B2(n401), .ZN(
        data_result[7]) );
  OAI22_X1 U860 ( .A1(n375), .A2(n611), .B1(n633), .B2(n402), .ZN(
        data_result[8]) );
  OAI22_X1 U861 ( .A1(n376), .A2(n634), .B1(n632), .B2(n403), .ZN(
        data_result[9]) );
  OAI22_X1 U862 ( .A1(n388), .A2(n634), .B1(n633), .B2(n405), .ZN(
        data_result[21]) );
  OAI22_X1 U863 ( .A1(n389), .A2(n634), .B1(n632), .B2(n406), .ZN(
        data_result[22]) );
  OAI22_X1 U864 ( .A1(n387), .A2(n634), .B1(n633), .B2(n404), .ZN(
        data_result[20]) );
  NAND4_X1 U865 ( .A1(n546), .A2(n547), .A3(n548), .A4(n549), .ZN(n523) );
  NOR4_X1 U866 ( .A1(n420), .A2(n421), .A3(n422), .A4(n423), .ZN(n546) );
  NOR4_X1 U867 ( .A1(n416), .A2(n417), .A3(n418), .A4(n419), .ZN(n547) );
  NOR4_X1 U868 ( .A1(n554), .A2(n555), .A3(n410), .A4(n411), .ZN(n548) );
  NAND4_X1 U869 ( .A1(n506), .A2(n505), .A3(n504), .A4(n503), .ZN(n534) );
  NAND4_X1 U870 ( .A1(n502), .A2(n501), .A3(n500), .A4(n499), .ZN(n533) );
  NAND4_X1 U871 ( .A1(n493), .A2(n492), .A3(n491), .A4(n490), .ZN(n532) );
  NAND4_X1 U872 ( .A1(n411), .A2(n412), .A3(n413), .A4(n414), .ZN(n542) );
  NAND4_X1 U873 ( .A1(n403), .A2(n404), .A3(n405), .A4(n406), .ZN(n531) );
  NAND4_X1 U874 ( .A1(n431), .A2(n432), .A3(n433), .A4(n434), .ZN(n544) );
  NAND4_X1 U875 ( .A1(n399), .A2(n400), .A3(n401), .A4(n402), .ZN(n528) );
  INV_X1 U876 ( .A(n509), .ZN(data_result[0]) );
  INV_X1 U877 ( .A(n490), .ZN(data_result[2]) );
  INV_X1 U878 ( .A(n499), .ZN(data_result[19]) );
  INV_X1 U879 ( .A(n503), .ZN(data_result[15]) );
  INV_X1 U880 ( .A(n504), .ZN(data_result[14]) );
  INV_X1 U881 ( .A(n500), .ZN(data_result[18]) );
  INV_X1 U882 ( .A(n491), .ZN(data_result[29]) );
  INV_X1 U883 ( .A(n505), .ZN(data_result[13]) );
  INV_X1 U884 ( .A(n501), .ZN(data_result[17]) );
  INV_X1 U885 ( .A(n492), .ZN(data_result[28]) );
  INV_X1 U886 ( .A(n498), .ZN(data_result[1]) );
  INV_X1 U887 ( .A(n506), .ZN(data_result[12]) );
  INV_X1 U888 ( .A(n502), .ZN(data_result[16]) );
  INV_X1 U889 ( .A(n493), .ZN(data_result[27]) );
  INV_X1 U890 ( .A(n507), .ZN(data_result[11]) );
  INV_X1 U891 ( .A(n508), .ZN(data_result[10]) );
  OAI22_X1 U892 ( .A1(data_operandA[4]), .A2(n675), .B1(product_out[5]), .B2(
        n673), .ZN(n583) );
  OAI22_X1 U893 ( .A1(data_operandA[5]), .A2(n675), .B1(product_out[6]), .B2(
        n673), .ZN(n584) );
  OAI22_X1 U894 ( .A1(data_operandA[8]), .A2(n675), .B1(product_out[9]), .B2(
        n672), .ZN(n587) );
  OAI22_X1 U895 ( .A1(data_operandA[2]), .A2(n675), .B1(product_out[3]), .B2(
        n673), .ZN(n581) );
  OAI22_X1 U896 ( .A1(data_operandA[7]), .A2(n675), .B1(product_out[8]), .B2(
        n672), .ZN(n586) );
  OAI22_X1 U897 ( .A1(data_operandA[3]), .A2(n675), .B1(product_out[4]), .B2(
        n673), .ZN(n582) );
  OAI22_X1 U898 ( .A1(data_operandA[6]), .A2(n675), .B1(product_out[7]), .B2(
        n672), .ZN(n585) );
  INV_X1 U899 ( .A(n478), .ZN(n390) );
  AOI22_X1 U900 ( .A1(data_operandA[31]), .A2(sign_fixed[23]), .B1(n681), .B2(
        data_operandA[23]), .ZN(n478) );
  AOI22_X1 U901 ( .A1(n649), .A2(data_operandB[12]), .B1(n668), .B2(
        data_operandA[12]), .ZN(n575) );
  AOI22_X1 U902 ( .A1(n649), .A2(data_operandB[10]), .B1(n668), .B2(
        data_operandA[10]), .ZN(n577) );
  INV_X1 U903 ( .A(n483), .ZN(n395) );
  AOI22_X1 U904 ( .A1(data_operandA[31]), .A2(sign_fixed[28]), .B1(n681), .B2(
        data_operandA[28]), .ZN(n483) );
  INV_X1 U905 ( .A(n481), .ZN(n393) );
  AOI22_X1 U906 ( .A1(data_operandA[31]), .A2(sign_fixed[26]), .B1(n681), .B2(
        data_operandA[26]), .ZN(n481) );
  INV_X1 U907 ( .A(n479), .ZN(n391) );
  AOI22_X1 U908 ( .A1(data_operandA[31]), .A2(sign_fixed[24]), .B1(n681), .B2(
        data_operandA[24]), .ZN(n479) );
  AOI22_X1 U909 ( .A1(n649), .A2(data_operandB[1]), .B1(n645), .B2(
        data_operandA[1]), .ZN(n567) );
  BUF_X1 U910 ( .A(ctrl_DIV), .Z(n672) );
  INV_X1 U911 ( .A(product_out[35]), .ZN(n410) );
  INV_X1 U912 ( .A(product_out[36]), .ZN(n411) );
  INV_X1 U913 ( .A(sign_fixed[31]), .ZN(n398) );
  INV_X1 U914 ( .A(product_out[34]), .ZN(n409) );
  INV_X1 U915 ( .A(product_out[33]), .ZN(n408) );
  INV_X1 U916 ( .A(product_out[32]), .ZN(n407) );
  INV_X1 U917 ( .A(data_operandB[5]), .ZN(n458) );
  INV_X1 U918 ( .A(data_operandB[7]), .ZN(n456) );
  INV_X1 U919 ( .A(data_operandA[5]), .ZN(n448) );
  INV_X1 U920 ( .A(data_operandA[6]), .ZN(n447) );
  INV_X1 U921 ( .A(data_operandA[7]), .ZN(n446) );
  INV_X1 U922 ( .A(data_operandB[6]), .ZN(n457) );
  INV_X1 U923 ( .A(n484), .ZN(n396) );
  AOI22_X1 U924 ( .A1(data_operandA[31]), .A2(sign_fixed[29]), .B1(n681), .B2(
        data_operandA[29]), .ZN(n484) );
  INV_X1 U925 ( .A(n482), .ZN(n394) );
  AOI22_X1 U926 ( .A1(data_operandA[31]), .A2(sign_fixed[27]), .B1(n681), .B2(
        data_operandA[27]), .ZN(n482) );
  INV_X1 U927 ( .A(n480), .ZN(n392) );
  AOI22_X1 U928 ( .A1(data_operandA[31]), .A2(sign_fixed[25]), .B1(n681), .B2(
        data_operandA[25]), .ZN(n480) );
  OAI22_X1 U929 ( .A1(data_operandA[26]), .A2(n677), .B1(product_out[27]), 
        .B2(n669), .ZN(n605) );
  OAI22_X1 U930 ( .A1(data_operandA[24]), .A2(n677), .B1(product_out[25]), 
        .B2(n669), .ZN(n603) );
  OAI22_X1 U931 ( .A1(data_operandA[13]), .A2(n676), .B1(product_out[14]), 
        .B2(n671), .ZN(n592) );
  OAI22_X1 U932 ( .A1(data_operandA[21]), .A2(n676), .B1(product_out[22]), 
        .B2(n670), .ZN(n600) );
  OAI22_X1 U933 ( .A1(data_operandA[16]), .A2(n676), .B1(product_out[17]), 
        .B2(n671), .ZN(n595) );
  OAI22_X1 U934 ( .A1(data_operandA[20]), .A2(n676), .B1(product_out[21]), 
        .B2(n670), .ZN(n599) );
  OAI22_X1 U935 ( .A1(data_operandA[12]), .A2(n676), .B1(product_out[13]), 
        .B2(n671), .ZN(n591) );
  OAI22_X1 U936 ( .A1(data_operandA[10]), .A2(n675), .B1(product_out[11]), 
        .B2(n672), .ZN(n589) );
  OAI22_X1 U937 ( .A1(data_operandA[18]), .A2(n676), .B1(product_out[19]), 
        .B2(n670), .ZN(n597) );
  OAI22_X1 U938 ( .A1(data_operandA[29]), .A2(n677), .B1(product_out[30]), 
        .B2(n669), .ZN(n608) );
  OAI22_X1 U939 ( .A1(data_operandA[28]), .A2(n677), .B1(product_out[29]), 
        .B2(n669), .ZN(n607) );
  OAI22_X1 U940 ( .A1(data_operandA[23]), .A2(n676), .B1(product_out[24]), 
        .B2(n669), .ZN(n602) );
  OAI22_X1 U941 ( .A1(data_operandA[15]), .A2(n676), .B1(product_out[16]), 
        .B2(n671), .ZN(n594) );
  OAI22_X1 U942 ( .A1(data_operandA[31]), .A2(n677), .B1(product_out[32]), 
        .B2(n669), .ZN(n610) );
  OAI22_X1 U943 ( .A1(data_operandA[25]), .A2(n677), .B1(product_out[26]), 
        .B2(n669), .ZN(n604) );
  OAI22_X1 U944 ( .A1(data_operandA[30]), .A2(n677), .B1(product_out[31]), 
        .B2(n671), .ZN(n609) );
  OAI22_X1 U945 ( .A1(data_operandA[14]), .A2(n676), .B1(product_out[15]), 
        .B2(n671), .ZN(n593) );
  OAI22_X1 U946 ( .A1(data_operandA[11]), .A2(n675), .B1(product_out[12]), 
        .B2(n672), .ZN(n590) );
  OAI22_X1 U947 ( .A1(data_operandA[17]), .A2(n676), .B1(product_out[18]), 
        .B2(n670), .ZN(n596) );
  OAI22_X1 U948 ( .A1(data_operandA[19]), .A2(n676), .B1(product_out[20]), 
        .B2(n670), .ZN(n598) );
  OAI22_X1 U949 ( .A1(data_operandA[27]), .A2(n677), .B1(product_out[28]), 
        .B2(n669), .ZN(n606) );
  OAI22_X1 U950 ( .A1(data_operandA[9]), .A2(n675), .B1(product_out[10]), .B2(
        n672), .ZN(n588) );
  OAI22_X1 U951 ( .A1(data_operandA[22]), .A2(n676), .B1(product_out[23]), 
        .B2(n670), .ZN(n601) );
  BUF_X1 U952 ( .A(ctrl_DIV), .Z(n669) );
  BUF_X1 U953 ( .A(ctrl_DIV), .Z(n671) );
  AOI22_X1 U954 ( .A1(n649), .A2(data_operandB[19]), .B1(n661), .B2(
        data_operandA[19]), .ZN(n568) );
  AOI22_X1 U955 ( .A1(n618), .A2(data_operandB[28]), .B1(n662), .B2(
        data_operandA[28]), .ZN(n561) );
  AOI22_X1 U956 ( .A1(n648), .A2(data_operandB[16]), .B1(n667), .B2(
        data_operandA[16]), .ZN(n571) );
  AOI22_X1 U957 ( .A1(n648), .A2(data_operandB[29]), .B1(n664), .B2(
        data_operandA[29]), .ZN(n560) );
  AOI22_X1 U958 ( .A1(n649), .A2(data_operandB[18]), .B1(n662), .B2(
        data_operandA[18]), .ZN(n569) );
  INV_X1 U959 ( .A(n477), .ZN(n386) );
  AOI22_X1 U960 ( .A1(data_operandA[31]), .A2(sign_fixed[19]), .B1(n681), .B2(
        data_operandA[19]), .ZN(n477) );
  INV_X1 U961 ( .A(n476), .ZN(n385) );
  AOI22_X1 U962 ( .A1(data_operandA[31]), .A2(sign_fixed[18]), .B1(n681), .B2(
        data_operandA[18]), .ZN(n476) );
  INV_X1 U963 ( .A(n475), .ZN(n384) );
  AOI22_X1 U964 ( .A1(data_operandA[31]), .A2(sign_fixed[17]), .B1(n681), .B2(
        data_operandA[17]), .ZN(n475) );
  AOI22_X1 U965 ( .A1(n618), .A2(data_operandB[25]), .B1(n664), .B2(
        data_operandA[25]), .ZN(n564) );
  AOI22_X1 U966 ( .A1(n648), .A2(data_operandB[27]), .B1(n664), .B2(
        data_operandA[27]), .ZN(n562) );
  INV_X1 U967 ( .A(n466), .ZN(n370) );
  AOI22_X1 U968 ( .A1(data_operandA[31]), .A2(sign_fixed[3]), .B1(n681), .B2(
        data_operandA[3]), .ZN(n466) );
  BUF_X1 U969 ( .A(ctrl_DIV), .Z(n670) );
  INV_X1 U970 ( .A(product_out[47]), .ZN(n422) );
  INV_X1 U971 ( .A(product_out[43]), .ZN(n418) );
  INV_X1 U972 ( .A(product_out[42]), .ZN(n417) );
  INV_X1 U973 ( .A(product_out[46]), .ZN(n421) );
  INV_X1 U974 ( .A(product_out[41]), .ZN(n416) );
  INV_X1 U975 ( .A(product_out[45]), .ZN(n420) );
  INV_X1 U976 ( .A(product_out[44]), .ZN(n419) );
  INV_X1 U977 ( .A(sign_fixed[20]), .ZN(n387) );
  INV_X1 U978 ( .A(product_out[39]), .ZN(n414) );
  INV_X1 U979 ( .A(product_out[59]), .ZN(n434) );
  INV_X1 U980 ( .A(product_out[48]), .ZN(n423) );
  INV_X1 U981 ( .A(product_out[38]), .ZN(n413) );
  INV_X1 U982 ( .A(product_out[58]), .ZN(n433) );
  INV_X1 U983 ( .A(product_out[37]), .ZN(n412) );
  INV_X1 U984 ( .A(product_out[57]), .ZN(n432) );
  INV_X1 U985 ( .A(product_out[40]), .ZN(n415) );
  INV_X1 U986 ( .A(product_out[56]), .ZN(n431) );
  INV_X1 U987 ( .A(product_out[63]), .ZN(n438) );
  INV_X1 U988 ( .A(product_out[62]), .ZN(n437) );
  INV_X1 U989 ( .A(product_out[53]), .ZN(n428) );
  INV_X1 U990 ( .A(product_out[49]), .ZN(n424) );
  INV_X1 U991 ( .A(product_out[61]), .ZN(n436) );
  INV_X1 U992 ( .A(product_out[50]), .ZN(n425) );
  INV_X1 U993 ( .A(product_out[54]), .ZN(n429) );
  INV_X1 U994 ( .A(product_out[51]), .ZN(n426) );
  INV_X1 U995 ( .A(product_out[55]), .ZN(n430) );
  INV_X1 U996 ( .A(product_out[52]), .ZN(n427) );
  INV_X1 U997 ( .A(product_out[60]), .ZN(n435) );
  INV_X1 U998 ( .A(sign_fixed[7]), .ZN(n374) );
  INV_X1 U999 ( .A(data_operandB[9]), .ZN(n454) );
  INV_X1 U1000 ( .A(sign_fixed[21]), .ZN(n388) );
  INV_X1 U1001 ( .A(sign_fixed[5]), .ZN(n372) );
  INV_X1 U1002 ( .A(sign_fixed[8]), .ZN(n375) );
  INV_X1 U1003 ( .A(data_operandB[8]), .ZN(n455) );
  INV_X1 U1004 ( .A(data_operandB[22]), .ZN(n451) );
  INV_X1 U1005 ( .A(data_operandB[21]), .ZN(n452) );
  INV_X1 U1006 ( .A(data_operandA[8]), .ZN(n445) );
  INV_X1 U1007 ( .A(data_operandA[9]), .ZN(n444) );
  INV_X1 U1008 ( .A(data_operandA[20]), .ZN(n443) );
  INV_X1 U1009 ( .A(data_operandA[21]), .ZN(n442) );
  INV_X1 U1010 ( .A(data_operandA[22]), .ZN(n441) );
  INV_X1 U1011 ( .A(data_operandB[20]), .ZN(n453) );
  INV_X1 U1012 ( .A(data_operandB[31]), .ZN(n449) );
  INV_X1 U1013 ( .A(product_out[64]), .ZN(n439) );
  INV_X1 U1014 ( .A(n474), .ZN(n383) );
  AOI22_X1 U1015 ( .A1(data_operandA[31]), .A2(sign_fixed[16]), .B1(n681), 
        .B2(data_operandA[16]), .ZN(n474) );
  INV_X1 U1016 ( .A(n469), .ZN(n378) );
  AOI22_X1 U1017 ( .A1(data_operandA[31]), .A2(sign_fixed[11]), .B1(n681), 
        .B2(data_operandA[11]), .ZN(n469) );
  INV_X1 U1018 ( .A(n468), .ZN(n377) );
  AOI22_X1 U1019 ( .A1(data_operandA[31]), .A2(sign_fixed[10]), .B1(n681), 
        .B2(data_operandA[10]), .ZN(n468) );
  INV_X1 U1020 ( .A(n473), .ZN(n382) );
  AOI22_X1 U1021 ( .A1(data_operandA[31]), .A2(sign_fixed[15]), .B1(n681), 
        .B2(data_operandA[15]), .ZN(n473) );
  INV_X1 U1022 ( .A(n472), .ZN(n381) );
  AOI22_X1 U1023 ( .A1(data_operandA[31]), .A2(sign_fixed[14]), .B1(n681), 
        .B2(data_operandA[14]), .ZN(n472) );
  INV_X1 U1024 ( .A(n471), .ZN(n380) );
  AOI22_X1 U1025 ( .A1(data_operandA[31]), .A2(sign_fixed[13]), .B1(n681), 
        .B2(data_operandA[13]), .ZN(n471) );
  INV_X1 U1026 ( .A(n470), .ZN(n379) );
  AOI22_X1 U1027 ( .A1(data_operandA[31]), .A2(sign_fixed[12]), .B1(n681), 
        .B2(data_operandA[12]), .ZN(n470) );
  INV_X1 U1028 ( .A(n467), .ZN(n371) );
  AOI22_X1 U1029 ( .A1(data_operandA[31]), .A2(sign_fixed[4]), .B1(n681), .B2(
        data_operandA[4]), .ZN(n467) );
  INV_X1 U1030 ( .A(n465), .ZN(n369) );
  AOI22_X1 U1031 ( .A1(data_operandA[31]), .A2(sign_fixed[2]), .B1(n680), .B2(
        data_operandA[2]), .ZN(n465) );
  INV_X1 U1032 ( .A(n464), .ZN(n368) );
  AOI22_X1 U1033 ( .A1(data_operandA[31]), .A2(sign_fixed[1]), .B1(n680), .B2(
        data_operandA[1]), .ZN(n464) );
  INV_X1 U1034 ( .A(n463), .ZN(n367) );
  AOI22_X1 U1035 ( .A1(data_operandA[31]), .A2(sign_fixed[0]), .B1(n680), .B2(
        data_operandA[0]), .ZN(n463) );
  INV_X1 U1036 ( .A(op_div), .ZN(n340) );
  NOR4_X1 U1037 ( .A1(n550), .A2(n551), .A3(n552), .A4(n553), .ZN(n549) );
  NAND4_X1 U1038 ( .A1(product_out[56]), .A2(product_out[55]), .A3(
        product_out[54]), .A4(product_out[53]), .ZN(n551) );
  NAND4_X1 U1039 ( .A1(product_out[64]), .A2(product_out[63]), .A3(
        product_out[62]), .A4(product_out[61]), .ZN(n553) );
  NAND4_X1 U1040 ( .A1(product_out[52]), .A2(product_out[51]), .A3(
        product_out[50]), .A4(product_out[49]), .ZN(n550) );
  NOR4_X1 U1041 ( .A1(n514), .A2(n515), .A3(n516), .A4(n517), .ZN(n513) );
  OR4_X1 U1042 ( .A1(data_operandB[28]), .A2(data_operandB[29]), .A3(
        data_operandB[2]), .A4(data_operandB[30]), .ZN(n516) );
  OR4_X1 U1043 ( .A1(data_operandB[24]), .A2(data_operandB[25]), .A3(
        data_operandB[26]), .A4(data_operandB[27]), .ZN(n517) );
  NAND4_X1 U1044 ( .A1(n457), .A2(n456), .A3(n455), .A4(n454), .ZN(n514) );
  NOR4_X1 U1045 ( .A1(n518), .A2(n519), .A3(n520), .A4(n521), .ZN(n512) );
  OR4_X1 U1046 ( .A1(data_operandB[17]), .A2(data_operandB[18]), .A3(
        data_operandB[19]), .A4(data_operandB[1]), .ZN(n519) );
  OR4_X1 U1047 ( .A1(data_operandB[13]), .A2(data_operandB[14]), .A3(
        data_operandB[15]), .A4(data_operandB[16]), .ZN(n520) );
  OR4_X1 U1048 ( .A1(data_operandB[0]), .A2(data_operandB[10]), .A3(
        data_operandB[11]), .A4(data_operandB[12]), .ZN(n521) );
  AOI22_X1 U1049 ( .A1(sign_fixed[19]), .A2(n633), .B1(n634), .B2(
        product_out[20]), .ZN(n499) );
  AOI22_X1 U1050 ( .A1(sign_fixed[2]), .A2(n633), .B1(n611), .B2(
        product_out[3]), .ZN(n490) );
  AOI22_X1 U1051 ( .A1(sign_fixed[15]), .A2(n632), .B1(n634), .B2(
        product_out[16]), .ZN(n503) );
  AOI22_X1 U1052 ( .A1(sign_fixed[14]), .A2(n633), .B1(n611), .B2(
        product_out[15]), .ZN(n504) );
  AOI22_X1 U1053 ( .A1(sign_fixed[18]), .A2(n633), .B1(n634), .B2(
        product_out[19]), .ZN(n500) );
  AOI22_X1 U1054 ( .A1(sign_fixed[29]), .A2(n633), .B1(n611), .B2(
        product_out[30]), .ZN(n491) );
  AOI22_X1 U1055 ( .A1(sign_fixed[13]), .A2(n633), .B1(n611), .B2(
        product_out[14]), .ZN(n505) );
  AOI22_X1 U1056 ( .A1(sign_fixed[17]), .A2(n633), .B1(n634), .B2(
        product_out[18]), .ZN(n501) );
  AOI22_X1 U1057 ( .A1(sign_fixed[28]), .A2(n633), .B1(n611), .B2(
        product_out[29]), .ZN(n492) );
  AOI22_X1 U1058 ( .A1(sign_fixed[12]), .A2(n633), .B1(n611), .B2(
        product_out[13]), .ZN(n506) );
  AOI22_X1 U1059 ( .A1(sign_fixed[16]), .A2(n633), .B1(n634), .B2(
        product_out[17]), .ZN(n502) );
  AOI22_X1 U1060 ( .A1(sign_fixed[27]), .A2(n633), .B1(n611), .B2(
        product_out[28]), .ZN(n493) );
  AOI22_X1 U1061 ( .A1(sign_fixed[11]), .A2(n632), .B1(n634), .B2(
        product_out[12]), .ZN(n507) );
  AOI22_X1 U1062 ( .A1(sign_fixed[10]), .A2(n632), .B1(n611), .B2(
        product_out[11]), .ZN(n508) );
  OAI22_X1 U1063 ( .A1(div_ready), .A2(n510), .B1(n511), .B2(n339), .ZN(
        data_exception) );
  AOI21_X1 U1064 ( .B1(n512), .B2(n513), .A(div_sign_ovf), .ZN(n511) );
  AOI221_X1 U1065 ( .B1(n522), .B2(data_result[31]), .C1(n523), .C2(n524), .A(
        n525), .ZN(n510) );
  NAND4_X1 U1066 ( .A1(n536), .A2(n537), .A3(n538), .A4(n539), .ZN(n524) );
  NOR4_X1 U1067 ( .A1(product_out[51]), .A2(product_out[50]), .A3(
        product_out[49]), .A4(product_out[48]), .ZN(n536) );
  NOR4_X1 U1068 ( .A1(product_out[55]), .A2(product_out[54]), .A3(
        product_out[53]), .A4(product_out[52]), .ZN(n537) );
  NOR4_X1 U1069 ( .A1(n544), .A2(n545), .A3(product_out[61]), .A4(
        product_out[60]), .ZN(n538) );
  NAND4_X1 U1070 ( .A1(product_out[60]), .A2(product_out[59]), .A3(
        product_out[58]), .A4(product_out[57]), .ZN(n552) );
  NAND4_X1 U1071 ( .A1(product_out[40]), .A2(product_out[39]), .A3(
        product_out[38]), .A4(product_out[37]), .ZN(n554) );
  NAND4_X1 U1072 ( .A1(n449), .A2(n460), .A3(n459), .A4(n458), .ZN(n515) );
  INV_X1 U1073 ( .A(data_operandB[3]), .ZN(n460) );
  INV_X1 U1074 ( .A(data_operandB[4]), .ZN(n459) );
  NAND4_X1 U1075 ( .A1(n453), .A2(n452), .A3(n451), .A4(n450), .ZN(n518) );
  INV_X1 U1076 ( .A(data_operandB[23]), .ZN(n450) );
  OR4_X1 U1077 ( .A1(product_out[24]), .A2(product_out[25]), .A3(
        product_out[26]), .A4(product_out[27]), .ZN(n530) );
  INV_X1 U1078 ( .A(product_out[23]), .ZN(n406) );
  INV_X1 U1079 ( .A(product_out[9]), .ZN(n402) );
  INV_X1 U1080 ( .A(product_out[22]), .ZN(n405) );
  INV_X1 U1081 ( .A(product_out[8]), .ZN(n401) );
  INV_X1 U1082 ( .A(product_out[21]), .ZN(n404) );
  INV_X1 U1083 ( .A(product_out[7]), .ZN(n400) );
  INV_X1 U1084 ( .A(product_out[10]), .ZN(n403) );
  INV_X1 U1085 ( .A(product_out[6]), .ZN(n399) );
  INV_X1 U1086 ( .A(div_ready), .ZN(n339) );
  INV_X1 U1087 ( .A(n494), .ZN(data_result[26]) );
  AOI22_X1 U1088 ( .A1(sign_fixed[26]), .A2(n632), .B1(n634), .B2(
        product_out[27]), .ZN(n494) );
  INV_X1 U1089 ( .A(n497), .ZN(data_result[23]) );
  AOI22_X1 U1090 ( .A1(sign_fixed[23]), .A2(n632), .B1(n611), .B2(
        product_out[24]), .ZN(n497) );
  INV_X1 U1091 ( .A(n496), .ZN(data_result[24]) );
  AOI22_X1 U1092 ( .A1(sign_fixed[24]), .A2(n632), .B1(n634), .B2(
        product_out[25]), .ZN(n496) );
  INV_X1 U1093 ( .A(n495), .ZN(data_result[25]) );
  AOI22_X1 U1094 ( .A1(sign_fixed[25]), .A2(n632), .B1(n634), .B2(
        product_out[26]), .ZN(n495) );
  INV_X1 U1095 ( .A(n489), .ZN(data_result[30]) );
  AOI22_X1 U1096 ( .A1(sign_fixed[30]), .A2(n632), .B1(n634), .B2(
        product_out[31]), .ZN(n489) );
  INV_X1 U1097 ( .A(n488), .ZN(data_result[3]) );
  AOI22_X1 U1098 ( .A1(sign_fixed[3]), .A2(n632), .B1(n611), .B2(
        product_out[4]), .ZN(n488) );
  INV_X1 U1099 ( .A(n487), .ZN(data_result[4]) );
  AOI22_X1 U1100 ( .A1(sign_fixed[4]), .A2(n632), .B1(n634), .B2(
        product_out[5]), .ZN(n487) );
  BUF_X1 U1101 ( .A(n647), .Z(n644) );
  BUF_X1 U1102 ( .A(n646), .Z(n643) );
  INV_X1 U1103 ( .A(n621), .ZN(n652) );
  INV_X1 U1104 ( .A(n557), .ZN(n342) );
  AOI22_X1 U1105 ( .A1(n649), .A2(data_operandB[3]), .B1(n666), .B2(
        data_operandA[3]), .ZN(n557) );
  INV_X1 U1106 ( .A(n668), .ZN(n654) );
  AOI22_X1 U1107 ( .A1(sign_fixed[0]), .A2(n632), .B1(n611), .B2(n619), .ZN(
        n509) );
  INV_X1 U1108 ( .A(ctrl_MULT), .ZN(n461) );
  OR4_X1 U1109 ( .A1(n624), .A2(product_out[31]), .A3(product_out[4]), .A4(
        product_out[5]), .ZN(n529) );
  AOI22_X1 U1110 ( .A1(sign_fixed[1]), .A2(n632), .B1(n611), .B2(n624), .ZN(
        n498) );
  INV_X1 U1111 ( .A(n567), .ZN(n352) );
  INV_X1 U1112 ( .A(n578), .ZN(n363) );
  INV_X1 U1113 ( .A(n623), .ZN(n366) );
  AND2_X1 U1114 ( .A1(product_in[62]), .A2(n660), .ZN(n185) );
  AOI22_X1 U1115 ( .A1(n653), .A2(data_operandB[30]), .B1(n666), .B2(
        data_operandA[30]), .ZN(n558) );
  AOI22_X1 U1116 ( .A1(n653), .A2(data_operandB[26]), .B1(n664), .B2(
        data_operandA[26]), .ZN(n563) );
  AOI22_X1 U1117 ( .A1(n653), .A2(data_operandB[24]), .B1(n664), .B2(
        data_operandA[24]), .ZN(n565) );
  AOI22_X1 U1118 ( .A1(n653), .A2(data_operandB[23]), .B1(n664), .B2(
        data_operandA[23]), .ZN(n566) );
  AOI22_X1 U1119 ( .A1(n653), .A2(data_operandB[17]), .B1(n661), .B2(
        data_operandA[17]), .ZN(n570) );
  AOI22_X1 U1120 ( .A1(n653), .A2(data_operandB[15]), .B1(n667), .B2(
        data_operandA[15]), .ZN(n572) );
  AOI22_X1 U1121 ( .A1(n656), .A2(data_operandB[14]), .B1(n667), .B2(
        data_operandA[14]), .ZN(n573) );
  AOI22_X1 U1122 ( .A1(n655), .A2(data_operandB[13]), .B1(n667), .B2(
        data_operandA[13]), .ZN(n574) );
  AOI22_X1 U1123 ( .A1(n654), .A2(data_operandB[11]), .B1(n668), .B2(
        data_operandA[11]), .ZN(n576) );
  AOI22_X1 U1124 ( .A1(n648), .A2(data_operandB[4]), .B1(n666), .B2(
        data_operandA[4]), .ZN(n556) );
  AOI22_X1 U1125 ( .A1(n649), .A2(data_operandB[2]), .B1(n643), .B2(
        data_operandA[2]), .ZN(n559) );
  AOI22_X1 U1126 ( .A1(n652), .A2(data_operandB[0]), .B1(n645), .B2(
        data_operandA[0]), .ZN(n578) );
  INV_X2 U1127 ( .A(n668), .ZN(n653) );
  INV_X2 U1128 ( .A(n668), .ZN(n655) );
  INV_X1 U1129 ( .A(n621), .ZN(n648) );
  AOI22_X1 \ctrl/U24  ( .A1(div_ready), .A2(\ctrl/n18 ), .B1(\ctrl/mult_ready ), .B2(\ctrl/n17 ), .ZN(\ctrl/n8 ) );
  NOR3_X1 \ctrl/U23  ( .A1(\ctrl/decoded_seq[5] ), .A2(\ctrl/decoded_seq[4] ), 
        .A3(\ctrl/decoded_seq[6] ), .ZN(\ctrl/n10 ) );
  OAI21_X1 \ctrl/U22  ( .B1(\ctrl/decoded_seq[3] ), .B2(\ctrl/n14 ), .A(
        \ctrl/n22 ), .ZN(\ctrl/n7 ) );
  NOR2_X1 \ctrl/U21  ( .A1(n614), .A2(n615), .ZN(\ctrl/n11 ) );
  OR3_X1 \ctrl/U20  ( .A1(n615), .A2(\ctrl/decoded_seq[3] ), .A3(
        \ctrl/decoded_seq[2] ), .ZN(\ctrl/n12 ) );
  CLKBUF_X1 \ctrl/U18  ( .A(\ctrl/op_mult_int ), .Z(\ctrl/n22 ) );
  OR3_X1 \ctrl/U17  ( .A1(\ctrl/n15 ), .A2(\ctrl/n13 ), .A3(
        \ctrl/decoded_seq[4] ), .ZN(\ctrl/n20 ) );
  INV_X1 \ctrl/U16  ( .A(\ctrl/n22 ), .ZN(\ctrl/n19 ) );
  AND2_X1 \ctrl/U15  ( .A1(\ctrl/op_div_int ), .A2(\ctrl/n11 ), .ZN(op_div) );
  INV_X1 \ctrl/U14  ( .A(\ctrl/n8 ), .ZN(data_resultRDY) );
  NAND2_X1 \ctrl/U13  ( .A1(\ctrl/n11 ), .A2(\ctrl/n8 ), .ZN(\ctrl/n_3_net_ )
         );
  CLKBUF_X1 \ctrl/U12  ( .A(op_mult), .Z(\ctrl/n17 ) );
  INV_X1 \ctrl/U11  ( .A(\ctrl/n17 ), .ZN(\ctrl/n18 ) );
  CLKBUF_X1 \ctrl/U10  ( .A(\ctrl/decoded_seq[5] ), .Z(\ctrl/n15 ) );
  OR2_X1 \ctrl/U9  ( .A1(n614), .A2(n615), .ZN(\ctrl/n21 ) );
  OAI22_X1 \ctrl/U8  ( .A1(\ctrl/n22 ), .A2(\ctrl/n9 ), .B1(\ctrl/n10 ), .B2(
        \ctrl/n19 ), .ZN(operandA_shift_0_) );
  BUF_X1 \ctrl/U7  ( .A(\ctrl/decoded_seq[4] ), .Z(\ctrl/n14 ) );
  INV_X2 \ctrl/U6  ( .A(\ctrl/n7 ), .ZN(shift) );
  CLKBUF_X1 \ctrl/U5  ( .A(\ctrl/decoded_seq[6] ), .Z(\ctrl/n13 ) );
  NOR4_X2 \ctrl/U4  ( .A1(\ctrl/n12 ), .A2(\ctrl/n20 ), .A3(
        \ctrl/decoded_seq[1] ), .A4(\ctrl/n19 ), .ZN(nop) );
  AND2_X1 \ctrl/U3  ( .A1(\ctrl/op_mult_int ), .A2(\ctrl/n11 ), .ZN(op_mult)
         );
  XOR2_X1 \ctrl/U19  ( .A(data_operandB[31]), .B(product_out[63]), .Z(
        \ctrl/n9 ) );
  INV_X1 \ctrl/decoder/U19  ( .A(product_out[2]), .ZN(\ctrl/decoder/n1 ) );
  NOR3_X1 \ctrl/decoder/U18  ( .A1(\ctrl/decoder/n11 ), .A2(\ctrl/decoder/n9 ), 
        .A3(\ctrl/decoder/n8 ), .ZN(\ctrl/decoded_seq[3] ) );
  NOR3_X1 \ctrl/decoder/U17  ( .A1(\ctrl/decoder/n11 ), .A2(\ctrl/decoder/n8 ), 
        .A3(\ctrl/decoder/n4 ), .ZN(\ctrl/decoded_seq[2] ) );
  NOR3_X1 \ctrl/decoder/U16  ( .A1(\ctrl/decoder/n9 ), .A2(\ctrl/decoder/n8 ), 
        .A3(\ctrl/decoder/n5 ), .ZN(\ctrl/decoded_seq[1] ) );
  NOR3_X1 \ctrl/decoder/U15  ( .A1(\ctrl/decoder/n10 ), .A2(\ctrl/decoder/n8 ), 
        .A3(\ctrl/decoder/n5 ), .ZN(\ctrl/SYNOPSYS_UNCONNECTED_2 ) );
  NOR3_X1 \ctrl/decoder/U14  ( .A1(\ctrl/decoder/n3 ), .A2(\ctrl/decoder/n1 ), 
        .A3(product_out[1]), .ZN(\ctrl/decoded_seq[5] ) );
  NOR3_X1 \ctrl/decoder/U13  ( .A1(\ctrl/decoder/n6 ), .A2(product_out[1]), 
        .A3(product_out[0]), .ZN(\ctrl/decoded_seq[4] ) );
  INV_X1 \ctrl/decoder/U12  ( .A(product_out[1]), .ZN(\ctrl/decoder/n2 ) );
  NOR3_X1 \ctrl/decoder/U11  ( .A1(\ctrl/decoder/n2 ), .A2(\ctrl/decoder/n1 ), 
        .A3(product_out[0]), .ZN(\ctrl/decoded_seq[6] ) );
  NOR3_X1 \ctrl/decoder/U10  ( .A1(\ctrl/decoder/n7 ), .A2(\ctrl/decoder/n9 ), 
        .A3(\ctrl/decoder/n11 ), .ZN(\ctrl/SYNOPSYS_UNCONNECTED_1 ) );
  INV_X1 \ctrl/decoder/U9  ( .A(product_out[0]), .ZN(\ctrl/decoder/n3 ) );
  INV_X1 \ctrl/decoder/U8  ( .A(\ctrl/decoder/n5 ), .ZN(\ctrl/decoder/n11 ) );
  CLKBUF_X1 \ctrl/decoder/U7  ( .A(\ctrl/decoder/n4 ), .Z(\ctrl/decoder/n10 )
         );
  INV_X1 \ctrl/decoder/U6  ( .A(\ctrl/decoder/n4 ), .ZN(\ctrl/decoder/n9 ) );
  CLKBUF_X1 \ctrl/decoder/U5  ( .A(product_out[2]), .Z(\ctrl/decoder/n8 ) );
  INV_X1 \ctrl/decoder/U4  ( .A(\ctrl/decoder/n8 ), .ZN(\ctrl/decoder/n7 ) );
  INV_X1 \ctrl/decoder/U3  ( .A(product_out[2]), .ZN(\ctrl/decoder/n6 ) );
  CLKBUF_X1 \ctrl/decoder/U2  ( .A(product_out[1]), .Z(\ctrl/decoder/n5 ) );
  CLKBUF_X1 \ctrl/decoder/U1  ( .A(product_out[0]), .Z(\ctrl/decoder/n4 ) );
  INV_X1 \ctrl/counter/U1  ( .A(clock), .ZN(\ctrl/counter/n1 ) );
  INV_X1 \ctrl/counter/tff_0/U2  ( .A(\ctrl/counter/tff_0/data ), .ZN(
        \ctrl/counter/w1 ) );
  XOR2_X1 \ctrl/counter/tff_0/U3  ( .A(1'b1), .B(\ctrl/counter/tff_0/data ), 
        .Z(\ctrl/counter/tff_0/d ) );
  INV_X1 \ctrl/counter/tff_0/dffe/U4  ( .A(\ctrl/n21 ), .ZN(
        \ctrl/counter/tff_0/dffe/n7 ) );
  NAND2_X1 \ctrl/counter/tff_0/dffe/U3  ( .A1(1'b1), .A2(
        \ctrl/counter/tff_0/d ), .ZN(\ctrl/counter/tff_0/dffe/n6 ) );
  OAI21_X1 \ctrl/counter/tff_0/dffe/U2  ( .B1(1'b1), .B2(
        \ctrl/counter/tff_0/dffe/n5 ), .A(\ctrl/counter/tff_0/dffe/n6 ), .ZN(
        \ctrl/counter/tff_0/dffe/n1 ) );
  DFFR_X1 \ctrl/counter/tff_0/dffe/q_reg  ( .D(\ctrl/counter/tff_0/dffe/n1 ), 
        .CK(\ctrl/counter/n1 ), .RN(\ctrl/counter/tff_0/dffe/n7 ), .Q(
        \ctrl/counter/tff_0/data ), .QN(\ctrl/counter/tff_0/dffe/n5 ) );
  INV_X1 \ctrl/counter/tff_1/U2  ( .A(\ctrl/counter/tff_1/data ), .ZN(
        \ctrl/counter/w2 ) );
  XOR2_X1 \ctrl/counter/tff_1/U3  ( .A(1'b1), .B(\ctrl/counter/tff_1/data ), 
        .Z(\ctrl/counter/tff_1/d ) );
  INV_X1 \ctrl/counter/tff_1/dffe/U4  ( .A(\ctrl/n21 ), .ZN(
        \ctrl/counter/tff_1/dffe/n7 ) );
  NAND2_X1 \ctrl/counter/tff_1/dffe/U3  ( .A1(1'b1), .A2(
        \ctrl/counter/tff_1/d ), .ZN(\ctrl/counter/tff_1/dffe/n6 ) );
  OAI21_X1 \ctrl/counter/tff_1/dffe/U2  ( .B1(1'b1), .B2(
        \ctrl/counter/tff_1/dffe/n5 ), .A(\ctrl/counter/tff_1/dffe/n6 ), .ZN(
        \ctrl/counter/tff_1/dffe/n1 ) );
  DFFR_X1 \ctrl/counter/tff_1/dffe/q_reg  ( .D(\ctrl/counter/tff_1/dffe/n1 ), 
        .CK(\ctrl/counter/w1 ), .RN(\ctrl/counter/tff_1/dffe/n7 ), .Q(
        \ctrl/counter/tff_1/data ), .QN(\ctrl/counter/tff_1/dffe/n5 ) );
  INV_X1 \ctrl/counter/tff_2/U2  ( .A(\ctrl/counter/tff_2/data ), .ZN(
        \ctrl/counter/w3 ) );
  XOR2_X1 \ctrl/counter/tff_2/U3  ( .A(1'b1), .B(\ctrl/counter/tff_2/data ), 
        .Z(\ctrl/counter/tff_2/d ) );
  INV_X1 \ctrl/counter/tff_2/dffe/U4  ( .A(\ctrl/n21 ), .ZN(
        \ctrl/counter/tff_2/dffe/n7 ) );
  NAND2_X1 \ctrl/counter/tff_2/dffe/U3  ( .A1(1'b1), .A2(
        \ctrl/counter/tff_2/d ), .ZN(\ctrl/counter/tff_2/dffe/n6 ) );
  OAI21_X1 \ctrl/counter/tff_2/dffe/U2  ( .B1(1'b1), .B2(
        \ctrl/counter/tff_2/dffe/n5 ), .A(\ctrl/counter/tff_2/dffe/n6 ), .ZN(
        \ctrl/counter/tff_2/dffe/n1 ) );
  DFFR_X1 \ctrl/counter/tff_2/dffe/q_reg  ( .D(\ctrl/counter/tff_2/dffe/n1 ), 
        .CK(\ctrl/counter/w2 ), .RN(\ctrl/counter/tff_2/dffe/n7 ), .Q(
        \ctrl/counter/tff_2/data ), .QN(\ctrl/counter/tff_2/dffe/n5 ) );
  INV_X1 \ctrl/counter/tff_3/U2  ( .A(\ctrl/counter/tff_3/data ), .ZN(
        \ctrl/counter/w4 ) );
  XOR2_X1 \ctrl/counter/tff_3/U3  ( .A(1'b1), .B(\ctrl/counter/tff_3/data ), 
        .Z(\ctrl/counter/tff_3/d ) );
  INV_X1 \ctrl/counter/tff_3/dffe/U4  ( .A(\ctrl/n21 ), .ZN(
        \ctrl/counter/tff_3/dffe/n7 ) );
  NAND2_X1 \ctrl/counter/tff_3/dffe/U3  ( .A1(1'b1), .A2(
        \ctrl/counter/tff_3/d ), .ZN(\ctrl/counter/tff_3/dffe/n6 ) );
  OAI21_X1 \ctrl/counter/tff_3/dffe/U2  ( .B1(1'b1), .B2(
        \ctrl/counter/tff_3/dffe/n5 ), .A(\ctrl/counter/tff_3/dffe/n6 ), .ZN(
        \ctrl/counter/tff_3/dffe/n1 ) );
  DFFR_X1 \ctrl/counter/tff_3/dffe/q_reg  ( .D(\ctrl/counter/tff_3/dffe/n1 ), 
        .CK(\ctrl/counter/w3 ), .RN(\ctrl/counter/tff_3/dffe/n7 ), .Q(
        \ctrl/counter/tff_3/data ), .QN(\ctrl/counter/tff_3/dffe/n5 ) );
  INV_X1 \ctrl/counter/tff_4/U2  ( .A(\ctrl/counter/w5 ), .ZN(
        \ctrl/counter/w6 ) );
  XOR2_X1 \ctrl/counter/tff_4/U3  ( .A(1'b1), .B(\ctrl/counter/w5 ), .Z(
        \ctrl/counter/tff_4/d ) );
  INV_X1 \ctrl/counter/tff_4/dffe/U4  ( .A(\ctrl/n21 ), .ZN(
        \ctrl/counter/tff_4/dffe/n7 ) );
  NAND2_X1 \ctrl/counter/tff_4/dffe/U3  ( .A1(1'b1), .A2(
        \ctrl/counter/tff_4/d ), .ZN(\ctrl/counter/tff_4/dffe/n6 ) );
  OAI21_X1 \ctrl/counter/tff_4/dffe/U2  ( .B1(1'b1), .B2(
        \ctrl/counter/tff_4/dffe/n5 ), .A(\ctrl/counter/tff_4/dffe/n6 ), .ZN(
        \ctrl/counter/tff_4/dffe/n1 ) );
  DFFR_X1 \ctrl/counter/tff_4/dffe/q_reg  ( .D(\ctrl/counter/tff_4/dffe/n1 ), 
        .CK(\ctrl/counter/w4 ), .RN(\ctrl/counter/tff_4/dffe/n7 ), .Q(
        \ctrl/counter/w5 ), .QN(\ctrl/counter/tff_4/dffe/n5 ) );
  INV_X1 \ctrl/counter/tff_5/U2  ( .A(\ctrl/counter/w7 ), .ZN(
        \ctrl/counter/tff_5/data_not ) );
  XOR2_X1 \ctrl/counter/tff_5/U3  ( .A(1'b1), .B(\ctrl/counter/w7 ), .Z(
        \ctrl/counter/tff_5/d ) );
  INV_X1 \ctrl/counter/tff_5/dffe/U4  ( .A(\ctrl/n21 ), .ZN(
        \ctrl/counter/tff_5/dffe/n7 ) );
  NAND2_X1 \ctrl/counter/tff_5/dffe/U3  ( .A1(1'b1), .A2(
        \ctrl/counter/tff_5/d ), .ZN(\ctrl/counter/tff_5/dffe/n6 ) );
  OAI21_X1 \ctrl/counter/tff_5/dffe/U2  ( .B1(1'b1), .B2(
        \ctrl/counter/tff_5/dffe/n5 ), .A(\ctrl/counter/tff_5/dffe/n6 ), .ZN(
        \ctrl/counter/tff_5/dffe/n1 ) );
  DFFR_X1 \ctrl/counter/tff_5/dffe/q_reg  ( .D(\ctrl/counter/tff_5/dffe/n1 ), 
        .CK(\ctrl/counter/w6 ), .RN(\ctrl/counter/tff_5/dffe/n7 ), .Q(
        \ctrl/counter/w7 ), .QN(\ctrl/counter/tff_5/dffe/n5 ) );
  INV_X1 \ctrl/counter/output16_dff/U4  ( .A(\ctrl/n21 ), .ZN(
        \ctrl/counter/output16_dff/n7 ) );
  NAND2_X1 \ctrl/counter/output16_dff/U3  ( .A1(1'b1), .A2(\ctrl/counter/w5 ), 
        .ZN(\ctrl/counter/output16_dff/n6 ) );
  OAI21_X1 \ctrl/counter/output16_dff/U2  ( .B1(1'b1), .B2(
        \ctrl/counter/output16_dff/n5 ), .A(\ctrl/counter/output16_dff/n6 ), 
        .ZN(\ctrl/counter/output16_dff/n1 ) );
  DFFR_X1 \ctrl/counter/output16_dff/q_reg  ( .D(
        \ctrl/counter/output16_dff/n1 ), .CK(clock), .RN(
        \ctrl/counter/output16_dff/n7 ), .Q(\ctrl/mult_ready ), .QN(
        \ctrl/counter/output16_dff/n5 ) );
  INV_X1 \ctrl/counter/output32_dff/U4  ( .A(\ctrl/n21 ), .ZN(
        \ctrl/counter/output32_dff/n7 ) );
  NAND2_X1 \ctrl/counter/output32_dff/U3  ( .A1(1'b1), .A2(\ctrl/counter/w7 ), 
        .ZN(\ctrl/counter/output32_dff/n6 ) );
  OAI21_X1 \ctrl/counter/output32_dff/U2  ( .B1(1'b1), .B2(
        \ctrl/counter/output32_dff/n5 ), .A(\ctrl/counter/output32_dff/n6 ), 
        .ZN(\ctrl/counter/output32_dff/n1 ) );
  DFFR_X1 \ctrl/counter/output32_dff/q_reg  ( .D(
        \ctrl/counter/output32_dff/n1 ), .CK(clock), .RN(
        \ctrl/counter/output32_dff/n7 ), .Q(div_ready), .QN(
        \ctrl/counter/output32_dff/n5 ) );
  NAND2_X1 \ctrl/cur_mult/U4  ( .A1(\ctrl/n_3_net_ ), .A2(n615), .ZN(
        \ctrl/cur_mult/n3 ) );
  OAI21_X1 \ctrl/cur_mult/U3  ( .B1(\ctrl/n_3_net_ ), .B2(\ctrl/cur_mult/n4 ), 
        .A(\ctrl/cur_mult/n3 ), .ZN(\ctrl/cur_mult/n1 ) );
  INV_X1 \ctrl/cur_mult/U2  ( .A(1'b0), .ZN(\ctrl/cur_mult/n2 ) );
  DFFR_X1 \ctrl/cur_mult/q_reg  ( .D(\ctrl/cur_mult/n1 ), .CK(clock), .RN(
        \ctrl/cur_mult/n2 ), .Q(\ctrl/op_mult_int ), .QN(\ctrl/cur_mult/n4 )
         );
  INV_X1 \ctrl/cur_div/U4  ( .A(1'b0), .ZN(\ctrl/cur_div/n7 ) );
  NAND2_X1 \ctrl/cur_div/U3  ( .A1(\ctrl/n_3_net_ ), .A2(n614), .ZN(
        \ctrl/cur_div/n6 ) );
  OAI21_X1 \ctrl/cur_div/U2  ( .B1(\ctrl/n_3_net_ ), .B2(\ctrl/cur_div/n5 ), 
        .A(\ctrl/cur_div/n6 ), .ZN(\ctrl/cur_div/n1 ) );
  DFFR_X1 \ctrl/cur_div/q_reg  ( .D(\ctrl/cur_div/n1 ), .CK(clock), .RN(
        \ctrl/cur_div/n7 ), .Q(\ctrl/op_div_int ), .QN(\ctrl/cur_div/n5 ) );
  INV_X1 \a_inv/U32  ( .A(n363), .ZN(data_operandA_not[0]) );
  INV_X1 \a_inv/U31  ( .A(n622), .ZN(data_operandA_not[1]) );
  INV_X1 \a_inv/U30  ( .A(n342), .ZN(data_operandA_not[3]) );
  INV_X1 \a_inv/U29  ( .A(n344), .ZN(data_operandA_not[2]) );
  INV_X1 \a_inv/U28  ( .A(n355), .ZN(data_operandA_not[17]) );
  INV_X1 \a_inv/U27  ( .A(n346), .ZN(data_operandA_not[28]) );
  INV_X1 \a_inv/U26  ( .A(n348), .ZN(data_operandA_not[26]) );
  INV_X1 \a_inv/U25  ( .A(n350), .ZN(data_operandA_not[24]) );
  INV_X1 \a_inv/U24  ( .A(n351), .ZN(data_operandA_not[23]) );
  INV_X1 \a_inv/U23  ( .A(n_1_net__31_), .ZN(data_operandA_not[31]) );
  INV_X1 \a_inv/U22  ( .A(n_1_net__22_), .ZN(data_operandA_not[22]) );
  INV_X1 \a_inv/U21  ( .A(n347), .ZN(data_operandA_not[27]) );
  INV_X1 \a_inv/U20  ( .A(n349), .ZN(data_operandA_not[25]) );
  INV_X1 \a_inv/U19  ( .A(n343), .ZN(data_operandA_not[30]) );
  INV_X1 \a_inv/U18  ( .A(n345), .ZN(data_operandA_not[29]) );
  INV_X1 \a_inv/U17  ( .A(n354), .ZN(data_operandA_not[18]) );
  INV_X1 \a_inv/U16  ( .A(n353), .ZN(data_operandA_not[19]) );
  INV_X1 \a_inv/U15  ( .A(n356), .ZN(data_operandA_not[16]) );
  INV_X1 \a_inv/U14  ( .A(n_1_net__21_), .ZN(data_operandA_not[21]) );
  INV_X1 \a_inv/U13  ( .A(n_1_net__20_), .ZN(data_operandA_not[20]) );
  INV_X1 \a_inv/U12  ( .A(n361), .ZN(data_operandA_not[11]) );
  INV_X1 \a_inv/U11  ( .A(n357), .ZN(data_operandA_not[15]) );
  INV_X1 \a_inv/U10  ( .A(n_1_net__8_), .ZN(data_operandA_not[8]) );
  INV_X1 \a_inv/U9  ( .A(n360), .ZN(data_operandA_not[12]) );
  INV_X1 \a_inv/U8  ( .A(n359), .ZN(data_operandA_not[13]) );
  INV_X1 \a_inv/U7  ( .A(n358), .ZN(data_operandA_not[14]) );
  INV_X1 \a_inv/U6  ( .A(n362), .ZN(data_operandA_not[10]) );
  INV_X1 \a_inv/U5  ( .A(n_1_net__7_), .ZN(data_operandA_not[7]) );
  INV_X1 \a_inv/U4  ( .A(n341), .ZN(data_operandA_not[4]) );
  INV_X1 \a_inv/U3  ( .A(n_1_net__9_), .ZN(data_operandA_not[9]) );
  INV_X1 \a_inv/U2  ( .A(n_1_net__6_), .ZN(data_operandA_not[6]) );
  INV_X1 \a_inv/U1  ( .A(n_1_net__5_), .ZN(data_operandA_not[5]) );
  INV_X1 \add_sub_mux/U76  ( .A(\add_sub_mux/n65 ), .ZN(operandA[0]) );
  INV_X1 \add_sub_mux/U75  ( .A(\add_sub_mux/n54 ), .ZN(operandA[1]) );
  AOI22_X1 \add_sub_mux/U74  ( .A1(\add_sub_mux/n68 ), .A2(n626), .B1(
        \add_sub_mux/n70 ), .B2(data_operandA_not[0]), .ZN(\add_sub_mux/n65 )
         );
  AOI22_X1 \add_sub_mux/U73  ( .A1(\add_sub_mux/n66 ), .A2(n352), .B1(
        data_operandA_not[1]), .B2(\add_sub_mux/n75 ), .ZN(\add_sub_mux/n54 )
         );
  AOI22_X1 \add_sub_mux/U72  ( .A1(n342), .A2(\add_sub_mux/n72 ), .B1(
        data_operandA_not[3]), .B2(\add_sub_mux/n75 ), .ZN(\add_sub_mux/n40 )
         );
  AOI22_X1 \add_sub_mux/U71  ( .A1(n344), .A2(\add_sub_mux/n72 ), .B1(
        data_operandA_not[2]), .B2(\add_sub_mux/n75 ), .ZN(\add_sub_mux/n43 )
         );
  AOI22_X1 \add_sub_mux/U70  ( .A1(n362), .A2(\add_sub_mux/n67 ), .B1(
        data_operandA_not[10]), .B2(\add_sub_mux/n76 ), .ZN(\add_sub_mux/n64 )
         );
  AOI22_X1 \add_sub_mux/U69  ( .A1(n361), .A2(\add_sub_mux/n67 ), .B1(
        data_operandA_not[11]), .B2(\add_sub_mux/n69 ), .ZN(\add_sub_mux/n63 )
         );
  AOI22_X1 \add_sub_mux/U68  ( .A1(n360), .A2(\add_sub_mux/n67 ), .B1(
        data_operandA_not[12]), .B2(\add_sub_mux/n74 ), .ZN(\add_sub_mux/n62 )
         );
  AOI22_X1 \add_sub_mux/U67  ( .A1(n359), .A2(\add_sub_mux/n67 ), .B1(
        data_operandA_not[13]), .B2(\add_sub_mux/n74 ), .ZN(\add_sub_mux/n61 )
         );
  AOI22_X1 \add_sub_mux/U66  ( .A1(n358), .A2(\add_sub_mux/n67 ), .B1(
        data_operandA_not[14]), .B2(\add_sub_mux/n74 ), .ZN(\add_sub_mux/n60 )
         );
  AOI22_X1 \add_sub_mux/U65  ( .A1(n357), .A2(\add_sub_mux/n67 ), .B1(
        data_operandA_not[15]), .B2(\add_sub_mux/n76 ), .ZN(\add_sub_mux/n59 )
         );
  AOI22_X1 \add_sub_mux/U64  ( .A1(n356), .A2(\add_sub_mux/n67 ), .B1(
        data_operandA_not[16]), .B2(\add_sub_mux/n74 ), .ZN(\add_sub_mux/n58 )
         );
  AOI22_X1 \add_sub_mux/U63  ( .A1(n355), .A2(\add_sub_mux/n67 ), .B1(
        data_operandA_not[17]), .B2(\add_sub_mux/n76 ), .ZN(\add_sub_mux/n57 )
         );
  AOI22_X1 \add_sub_mux/U62  ( .A1(n354), .A2(\add_sub_mux/n67 ), .B1(
        data_operandA_not[18]), .B2(\add_sub_mux/n76 ), .ZN(\add_sub_mux/n56 )
         );
  AOI22_X1 \add_sub_mux/U61  ( .A1(n353), .A2(\add_sub_mux/n67 ), .B1(
        data_operandA_not[19]), .B2(\add_sub_mux/n74 ), .ZN(\add_sub_mux/n55 )
         );
  INV_X1 \add_sub_mux/U60  ( .A(\add_sub_mux/n40 ), .ZN(operandA[3]) );
  INV_X1 \add_sub_mux/U59  ( .A(\add_sub_mux/n57 ), .ZN(operandA[17]) );
  AOI22_X1 \add_sub_mux/U58  ( .A1(n346), .A2(\add_sub_mux/n71 ), .B1(
        data_operandA_not[28]), .B2(\add_sub_mux/n74 ), .ZN(\add_sub_mux/n45 )
         );
  INV_X1 \add_sub_mux/U57  ( .A(\add_sub_mux/n45 ), .ZN(operandA[28]) );
  AOI22_X1 \add_sub_mux/U56  ( .A1(n348), .A2(\add_sub_mux/n71 ), .B1(
        data_operandA_not[26]), .B2(\add_sub_mux/n74 ), .ZN(\add_sub_mux/n47 )
         );
  INV_X1 \add_sub_mux/U55  ( .A(\add_sub_mux/n47 ), .ZN(operandA[26]) );
  AOI22_X1 \add_sub_mux/U54  ( .A1(n350), .A2(\add_sub_mux/n71 ), .B1(
        data_operandA_not[24]), .B2(\add_sub_mux/n74 ), .ZN(\add_sub_mux/n49 )
         );
  INV_X1 \add_sub_mux/U53  ( .A(\add_sub_mux/n49 ), .ZN(operandA[24]) );
  AOI22_X1 \add_sub_mux/U52  ( .A1(n351), .A2(\add_sub_mux/n71 ), .B1(
        data_operandA_not[23]), .B2(\add_sub_mux/n74 ), .ZN(\add_sub_mux/n50 )
         );
  INV_X1 \add_sub_mux/U51  ( .A(\add_sub_mux/n50 ), .ZN(operandA[23]) );
  AOI22_X1 \add_sub_mux/U50  ( .A1(n_1_net__31_), .A2(\add_sub_mux/n71 ), .B1(
        data_operandA_not[31]), .B2(\add_sub_mux/n74 ), .ZN(\add_sub_mux/n41 )
         );
  INV_X1 \add_sub_mux/U49  ( .A(\add_sub_mux/n41 ), .ZN(operandA[31]) );
  AOI22_X1 \add_sub_mux/U48  ( .A1(n_1_net__22_), .A2(\add_sub_mux/n71 ), .B1(
        data_operandA_not[22]), .B2(\add_sub_mux/n74 ), .ZN(\add_sub_mux/n51 )
         );
  INV_X1 \add_sub_mux/U47  ( .A(\add_sub_mux/n51 ), .ZN(operandA[22]) );
  AOI22_X1 \add_sub_mux/U46  ( .A1(n347), .A2(\add_sub_mux/n71 ), .B1(
        data_operandA_not[27]), .B2(\add_sub_mux/n74 ), .ZN(\add_sub_mux/n46 )
         );
  INV_X1 \add_sub_mux/U45  ( .A(\add_sub_mux/n46 ), .ZN(operandA[27]) );
  AOI22_X1 \add_sub_mux/U44  ( .A1(n349), .A2(\add_sub_mux/n71 ), .B1(
        data_operandA_not[25]), .B2(\add_sub_mux/n74 ), .ZN(\add_sub_mux/n48 )
         );
  INV_X1 \add_sub_mux/U43  ( .A(\add_sub_mux/n48 ), .ZN(operandA[25]) );
  AOI22_X1 \add_sub_mux/U42  ( .A1(n343), .A2(\add_sub_mux/n71 ), .B1(
        data_operandA_not[30]), .B2(\add_sub_mux/n74 ), .ZN(\add_sub_mux/n42 )
         );
  INV_X1 \add_sub_mux/U41  ( .A(\add_sub_mux/n42 ), .ZN(operandA[30]) );
  AOI22_X1 \add_sub_mux/U40  ( .A1(n345), .A2(\add_sub_mux/n71 ), .B1(
        data_operandA_not[29]), .B2(\add_sub_mux/n74 ), .ZN(\add_sub_mux/n44 )
         );
  INV_X1 \add_sub_mux/U39  ( .A(\add_sub_mux/n44 ), .ZN(operandA[29]) );
  INV_X1 \add_sub_mux/U38  ( .A(\add_sub_mux/n56 ), .ZN(operandA[18]) );
  INV_X1 \add_sub_mux/U37  ( .A(\add_sub_mux/n55 ), .ZN(operandA[19]) );
  INV_X1 \add_sub_mux/U36  ( .A(\add_sub_mux/n58 ), .ZN(operandA[16]) );
  AOI22_X1 \add_sub_mux/U35  ( .A1(n_1_net__21_), .A2(\add_sub_mux/n71 ), .B1(
        data_operandA_not[21]), .B2(\add_sub_mux/n74 ), .ZN(\add_sub_mux/n52 )
         );
  INV_X1 \add_sub_mux/U34  ( .A(\add_sub_mux/n52 ), .ZN(operandA[21]) );
  AOI22_X1 \add_sub_mux/U33  ( .A1(n_1_net__20_), .A2(\add_sub_mux/n71 ), .B1(
        data_operandA_not[20]), .B2(\add_sub_mux/n74 ), .ZN(\add_sub_mux/n53 )
         );
  INV_X1 \add_sub_mux/U32  ( .A(\add_sub_mux/n53 ), .ZN(operandA[20]) );
  INV_X1 \add_sub_mux/U31  ( .A(\add_sub_mux/n63 ), .ZN(operandA[11]) );
  INV_X1 \add_sub_mux/U30  ( .A(\add_sub_mux/n59 ), .ZN(operandA[15]) );
  AOI22_X1 \add_sub_mux/U29  ( .A1(n_1_net__8_), .A2(\add_sub_mux/n71 ), .B1(
        data_operandA_not[8]), .B2(\add_sub_mux/n73 ), .ZN(\add_sub_mux/n35 )
         );
  INV_X1 \add_sub_mux/U28  ( .A(\add_sub_mux/n35 ), .ZN(operandA[8]) );
  INV_X1 \add_sub_mux/U27  ( .A(\add_sub_mux/n43 ), .ZN(operandA[2]) );
  INV_X1 \add_sub_mux/U26  ( .A(\add_sub_mux/n62 ), .ZN(operandA[12]) );
  INV_X1 \add_sub_mux/U25  ( .A(\add_sub_mux/n61 ), .ZN(operandA[13]) );
  INV_X1 \add_sub_mux/U24  ( .A(\add_sub_mux/n60 ), .ZN(operandA[14]) );
  INV_X1 \add_sub_mux/U23  ( .A(\add_sub_mux/n64 ), .ZN(operandA[10]) );
  AOI22_X1 \add_sub_mux/U22  ( .A1(n_1_net__7_), .A2(\add_sub_mux/n71 ), .B1(
        data_operandA_not[7]), .B2(\add_sub_mux/n73 ), .ZN(\add_sub_mux/n36 )
         );
  INV_X1 \add_sub_mux/U21  ( .A(\add_sub_mux/n36 ), .ZN(operandA[7]) );
  AOI22_X1 \add_sub_mux/U20  ( .A1(n341), .A2(\add_sub_mux/n33 ), .B1(
        data_operandA_not[4]), .B2(\add_sub_mux/n69 ), .ZN(\add_sub_mux/n39 )
         );
  INV_X1 \add_sub_mux/U19  ( .A(\add_sub_mux/n39 ), .ZN(operandA[4]) );
  AOI22_X1 \add_sub_mux/U18  ( .A1(n_1_net__9_), .A2(\add_sub_mux/n71 ), .B1(
        \add_sub_mux/n76 ), .B2(data_operandA_not[9]), .ZN(\add_sub_mux/n34 )
         );
  INV_X1 \add_sub_mux/U17  ( .A(\add_sub_mux/n34 ), .ZN(operandA[9]) );
  AOI22_X1 \add_sub_mux/U16  ( .A1(n_1_net__6_), .A2(\add_sub_mux/n71 ), .B1(
        data_operandA_not[6]), .B2(\add_sub_mux/n73 ), .ZN(\add_sub_mux/n37 )
         );
  INV_X1 \add_sub_mux/U15  ( .A(\add_sub_mux/n37 ), .ZN(operandA[6]) );
  AOI22_X1 \add_sub_mux/U14  ( .A1(n_1_net__5_), .A2(\add_sub_mux/n71 ), .B1(
        data_operandA_not[5]), .B2(\add_sub_mux/n73 ), .ZN(\add_sub_mux/n38 )
         );
  INV_X1 \add_sub_mux/U13  ( .A(\add_sub_mux/n38 ), .ZN(operandA[5]) );
  CLKBUF_X1 \add_sub_mux/U12  ( .A(\add_sub_mux/n69 ), .Z(\add_sub_mux/n73 )
         );
  BUF_X1 \add_sub_mux/U11  ( .A(operandA_shift_0_), .Z(\add_sub_mux/n70 ) );
  INV_X1 \add_sub_mux/U10  ( .A(\add_sub_mux/n70 ), .ZN(\add_sub_mux/n72 ) );
  INV_X1 \add_sub_mux/U9  ( .A(\add_sub_mux/n72 ), .ZN(\add_sub_mux/n69 ) );
  CLKBUF_X1 \add_sub_mux/U8  ( .A(\add_sub_mux/n69 ), .Z(\add_sub_mux/n76 ) );
  INV_X1 \add_sub_mux/U7  ( .A(operandA_shift_0_), .ZN(\add_sub_mux/n68 ) );
  INV_X1 \add_sub_mux/U6  ( .A(\add_sub_mux/n69 ), .ZN(\add_sub_mux/n67 ) );
  BUF_X1 \add_sub_mux/U5  ( .A(\add_sub_mux/n68 ), .Z(\add_sub_mux/n66 ) );
  INV_X1 \add_sub_mux/U4  ( .A(\add_sub_mux/n70 ), .ZN(\add_sub_mux/n71 ) );
  BUF_X1 \add_sub_mux/U3  ( .A(\add_sub_mux/n70 ), .Z(\add_sub_mux/n75 ) );
  CLKBUF_X1 \add_sub_mux/U2  ( .A(\add_sub_mux/n66 ), .Z(\add_sub_mux/n33 ) );
  CLKBUF_X2 \add_sub_mux/U1  ( .A(\add_sub_mux/n69 ), .Z(\add_sub_mux/n74 ) );
  AOI22_X1 \shift_booth_mux/U73  ( .A1(operandA[26]), .A2(
        \shift_booth_mux/n71 ), .B1(operandA[25]), .B2(\shift_booth_mux/n73 ), 
        .ZN(\shift_booth_mux/n90 ) );
  INV_X1 \shift_booth_mux/U72  ( .A(\shift_booth_mux/n90 ), .ZN(
        operandA_resolved[26]) );
  AOI22_X1 \shift_booth_mux/U71  ( .A1(operandA[27]), .A2(
        \shift_booth_mux/n71 ), .B1(operandA[26]), .B2(\shift_booth_mux/n73 ), 
        .ZN(\shift_booth_mux/n91 ) );
  INV_X1 \shift_booth_mux/U70  ( .A(\shift_booth_mux/n91 ), .ZN(
        operandA_resolved[27]) );
  AOI22_X1 \shift_booth_mux/U69  ( .A1(operandA[25]), .A2(
        \shift_booth_mux/n71 ), .B1(operandA[24]), .B2(\shift_booth_mux/n73 ), 
        .ZN(\shift_booth_mux/n89 ) );
  INV_X1 \shift_booth_mux/U68  ( .A(\shift_booth_mux/n89 ), .ZN(
        operandA_resolved[25]) );
  AOI22_X1 \shift_booth_mux/U67  ( .A1(operandA[24]), .A2(
        \shift_booth_mux/n71 ), .B1(operandA[23]), .B2(\shift_booth_mux/n73 ), 
        .ZN(\shift_booth_mux/n88 ) );
  INV_X1 \shift_booth_mux/U66  ( .A(\shift_booth_mux/n88 ), .ZN(
        operandA_resolved[24]) );
  AOI22_X1 \shift_booth_mux/U65  ( .A1(operandA[23]), .A2(
        \shift_booth_mux/n71 ), .B1(operandA[22]), .B2(\shift_booth_mux/n73 ), 
        .ZN(\shift_booth_mux/n87 ) );
  INV_X1 \shift_booth_mux/U64  ( .A(\shift_booth_mux/n87 ), .ZN(
        operandA_resolved[23]) );
  AOI22_X1 \shift_booth_mux/U63  ( .A1(operandA[31]), .A2(
        \shift_booth_mux/n71 ), .B1(operandA[30]), .B2(\shift_booth_mux/n73 ), 
        .ZN(\shift_booth_mux/n95 ) );
  INV_X1 \shift_booth_mux/U62  ( .A(\shift_booth_mux/n95 ), .ZN(
        operandA_resolved[31]) );
  AOI22_X1 \shift_booth_mux/U61  ( .A1(operandA[19]), .A2(
        \shift_booth_mux/n70 ), .B1(operandA[18]), .B2(\shift_booth_mux/n73 ), 
        .ZN(\shift_booth_mux/n83 ) );
  INV_X1 \shift_booth_mux/U60  ( .A(\shift_booth_mux/n83 ), .ZN(
        operandA_resolved[19]) );
  AOI22_X1 \shift_booth_mux/U59  ( .A1(operandA[22]), .A2(
        \shift_booth_mux/n71 ), .B1(operandA[21]), .B2(\shift_booth_mux/n73 ), 
        .ZN(\shift_booth_mux/n86 ) );
  INV_X1 \shift_booth_mux/U58  ( .A(\shift_booth_mux/n86 ), .ZN(
        operandA_resolved[22]) );
  AOI22_X1 \shift_booth_mux/U57  ( .A1(operandA[30]), .A2(
        \shift_booth_mux/n71 ), .B1(operandA[29]), .B2(\shift_booth_mux/n73 ), 
        .ZN(\shift_booth_mux/n94 ) );
  INV_X1 \shift_booth_mux/U56  ( .A(\shift_booth_mux/n94 ), .ZN(
        operandA_resolved[30]) );
  AOI22_X1 \shift_booth_mux/U55  ( .A1(operandA[16]), .A2(
        \shift_booth_mux/n70 ), .B1(operandA[15]), .B2(\shift_booth_mux/n73 ), 
        .ZN(\shift_booth_mux/n80 ) );
  INV_X1 \shift_booth_mux/U54  ( .A(\shift_booth_mux/n80 ), .ZN(
        operandA_resolved[16]) );
  AOI22_X1 \shift_booth_mux/U53  ( .A1(operandA[20]), .A2(
        \shift_booth_mux/n71 ), .B1(operandA[19]), .B2(\shift_booth_mux/n73 ), 
        .ZN(\shift_booth_mux/n84 ) );
  INV_X1 \shift_booth_mux/U52  ( .A(\shift_booth_mux/n84 ), .ZN(
        operandA_resolved[20]) );
  AOI22_X1 \shift_booth_mux/U51  ( .A1(operandA[21]), .A2(
        \shift_booth_mux/n71 ), .B1(operandA[20]), .B2(\shift_booth_mux/n73 ), 
        .ZN(\shift_booth_mux/n85 ) );
  INV_X1 \shift_booth_mux/U50  ( .A(\shift_booth_mux/n85 ), .ZN(
        operandA_resolved[21]) );
  AOI22_X1 \shift_booth_mux/U49  ( .A1(operandA[28]), .A2(
        \shift_booth_mux/n71 ), .B1(operandA[27]), .B2(\shift_booth_mux/n73 ), 
        .ZN(\shift_booth_mux/n92 ) );
  INV_X1 \shift_booth_mux/U48  ( .A(\shift_booth_mux/n92 ), .ZN(
        operandA_resolved[28]) );
  AOI22_X1 \shift_booth_mux/U47  ( .A1(operandA[29]), .A2(
        \shift_booth_mux/n71 ), .B1(operandA[28]), .B2(\shift_booth_mux/n73 ), 
        .ZN(\shift_booth_mux/n93 ) );
  INV_X1 \shift_booth_mux/U46  ( .A(\shift_booth_mux/n93 ), .ZN(
        operandA_resolved[29]) );
  AOI22_X1 \shift_booth_mux/U45  ( .A1(operandA[18]), .A2(
        \shift_booth_mux/n70 ), .B1(operandA[17]), .B2(\shift_booth_mux/n73 ), 
        .ZN(\shift_booth_mux/n82 ) );
  INV_X1 \shift_booth_mux/U44  ( .A(\shift_booth_mux/n82 ), .ZN(
        operandA_resolved[18]) );
  AOI22_X1 \shift_booth_mux/U43  ( .A1(operandA[17]), .A2(
        \shift_booth_mux/n70 ), .B1(operandA[16]), .B2(\shift_booth_mux/n73 ), 
        .ZN(\shift_booth_mux/n81 ) );
  INV_X1 \shift_booth_mux/U42  ( .A(\shift_booth_mux/n81 ), .ZN(
        operandA_resolved[17]) );
  AOI22_X1 \shift_booth_mux/U41  ( .A1(operandA[6]), .A2(\shift_booth_mux/n71 ), .B1(operandA[5]), .B2(\shift_booth_mux/n72 ), .ZN(\shift_booth_mux/n98 ) );
  INV_X1 \shift_booth_mux/U40  ( .A(\shift_booth_mux/n98 ), .ZN(
        operandA_resolved[6]) );
  AOI22_X1 \shift_booth_mux/U39  ( .A1(operandA[9]), .A2(\shift_booth_mux/n70 ), .B1(\shift_booth_mux/n69 ), .B2(operandA[8]), .ZN(\shift_booth_mux/n101 ) );
  INV_X1 \shift_booth_mux/U38  ( .A(\shift_booth_mux/n101 ), .ZN(
        operandA_resolved[9]) );
  AOI22_X1 \shift_booth_mux/U37  ( .A1(operandA[10]), .A2(
        \shift_booth_mux/n70 ), .B1(operandA[9]), .B2(\shift_booth_mux/n69 ), 
        .ZN(\shift_booth_mux/n74 ) );
  INV_X1 \shift_booth_mux/U36  ( .A(\shift_booth_mux/n74 ), .ZN(
        operandA_resolved[10]) );
  AOI22_X1 \shift_booth_mux/U35  ( .A1(operandA[12]), .A2(
        \shift_booth_mux/n70 ), .B1(operandA[11]), .B2(\shift_booth_mux/n73 ), 
        .ZN(\shift_booth_mux/n76 ) );
  INV_X1 \shift_booth_mux/U34  ( .A(\shift_booth_mux/n76 ), .ZN(
        operandA_resolved[12]) );
  AOI22_X1 \shift_booth_mux/U33  ( .A1(operandA[13]), .A2(
        \shift_booth_mux/n70 ), .B1(operandA[12]), .B2(\shift_booth_mux/n73 ), 
        .ZN(\shift_booth_mux/n77 ) );
  INV_X1 \shift_booth_mux/U32  ( .A(\shift_booth_mux/n77 ), .ZN(
        operandA_resolved[13]) );
  AOI22_X1 \shift_booth_mux/U31  ( .A1(operandA[15]), .A2(
        \shift_booth_mux/n70 ), .B1(operandA[14]), .B2(\shift_booth_mux/n73 ), 
        .ZN(\shift_booth_mux/n79 ) );
  INV_X1 \shift_booth_mux/U30  ( .A(\shift_booth_mux/n79 ), .ZN(
        operandA_resolved[15]) );
  AOI22_X1 \shift_booth_mux/U29  ( .A1(operandA[4]), .A2(\shift_booth_mux/n33 ), .B1(operandA[3]), .B2(\shift_booth_mux/n72 ), .ZN(\shift_booth_mux/n96 ) );
  INV_X1 \shift_booth_mux/U28  ( .A(\shift_booth_mux/n96 ), .ZN(
        operandA_resolved[4]) );
  AOI22_X1 \shift_booth_mux/U27  ( .A1(operandA[5]), .A2(\shift_booth_mux/n70 ), .B1(n612), .B2(\shift_booth_mux/n72 ), .ZN(\shift_booth_mux/n97 ) );
  INV_X1 \shift_booth_mux/U26  ( .A(\shift_booth_mux/n97 ), .ZN(
        operandA_resolved[5]) );
  AOI22_X1 \shift_booth_mux/U25  ( .A1(operandA[8]), .A2(\shift_booth_mux/n71 ), .B1(operandA[7]), .B2(\shift_booth_mux/n72 ), .ZN(\shift_booth_mux/n100 ) );
  INV_X1 \shift_booth_mux/U24  ( .A(\shift_booth_mux/n100 ), .ZN(
        operandA_resolved[8]) );
  AOI22_X1 \shift_booth_mux/U23  ( .A1(operandA[7]), .A2(\shift_booth_mux/n71 ), .B1(operandA[6]), .B2(\shift_booth_mux/n72 ), .ZN(\shift_booth_mux/n99 ) );
  INV_X1 \shift_booth_mux/U22  ( .A(\shift_booth_mux/n99 ), .ZN(
        operandA_resolved[7]) );
  AOI22_X1 \shift_booth_mux/U21  ( .A1(operandA[11]), .A2(
        \shift_booth_mux/n70 ), .B1(operandA[10]), .B2(\shift_booth_mux/n73 ), 
        .ZN(\shift_booth_mux/n75 ) );
  INV_X1 \shift_booth_mux/U20  ( .A(\shift_booth_mux/n75 ), .ZN(
        operandA_resolved[11]) );
  AOI22_X1 \shift_booth_mux/U19  ( .A1(operandA[14]), .A2(
        \shift_booth_mux/n70 ), .B1(operandA[13]), .B2(\shift_booth_mux/n73 ), 
        .ZN(\shift_booth_mux/n78 ) );
  INV_X1 \shift_booth_mux/U18  ( .A(\shift_booth_mux/n78 ), .ZN(
        operandA_resolved[14]) );
  INV_X1 \shift_booth_mux/U17  ( .A(\shift_booth_mux/n69 ), .ZN(
        \shift_booth_mux/n70 ) );
  INV_X1 \shift_booth_mux/U16  ( .A(\shift_booth_mux/n68 ), .ZN(
        \shift_booth_mux/n71 ) );
  MUX2_X1 \shift_booth_mux/U15  ( .A(operandA[2]), .B(operandA[1]), .S(shift), 
        .Z(operandA_resolved[2]) );
  NAND2_X1 \shift_booth_mux/U14  ( .A1(\shift_booth_mux/n66 ), .A2(
        \shift_booth_mux/n67 ), .ZN(operandA_resolved[1]) );
  NAND2_X1 \shift_booth_mux/U13  ( .A1(n627), .A2(shift), .ZN(
        \shift_booth_mux/n67 ) );
  NAND2_X1 \shift_booth_mux/U12  ( .A1(operandA[1]), .A2(\shift_booth_mux/n33 ), .ZN(\shift_booth_mux/n66 ) );
  NAND2_X1 \shift_booth_mux/U11  ( .A1(\shift_booth_mux/n54 ), .A2(
        \shift_booth_mux/n65 ), .ZN(operandA_resolved[0]) );
  NAND2_X1 \shift_booth_mux/U10  ( .A1(n629), .A2(shift), .ZN(
        \shift_booth_mux/n65 ) );
  NAND2_X1 \shift_booth_mux/U9  ( .A1(operandA[0]), .A2(\shift_booth_mux/n33 ), 
        .ZN(\shift_booth_mux/n54 ) );
  INV_X1 \shift_booth_mux/U8  ( .A(shift), .ZN(\shift_booth_mux/n33 ) );
  NAND2_X1 \shift_booth_mux/U7  ( .A1(\shift_booth_mux/n40 ), .A2(
        \shift_booth_mux/n43 ), .ZN(operandA_resolved[3]) );
  NAND2_X1 \shift_booth_mux/U6  ( .A1(n620), .A2(shift), .ZN(
        \shift_booth_mux/n43 ) );
  NAND2_X1 \shift_booth_mux/U5  ( .A1(operandA[3]), .A2(\shift_booth_mux/n33 ), 
        .ZN(\shift_booth_mux/n40 ) );
  CLKBUF_X1 \shift_booth_mux/U4  ( .A(shift), .Z(\shift_booth_mux/n68 ) );
  CLKBUF_X1 \shift_booth_mux/U3  ( .A(shift), .Z(\shift_booth_mux/n69 ) );
  BUF_X1 \shift_booth_mux/U2  ( .A(\shift_booth_mux/n68 ), .Z(
        \shift_booth_mux/n72 ) );
  CLKBUF_X3 \shift_booth_mux/U1  ( .A(\shift_booth_mux/n69 ), .Z(
        \shift_booth_mux/n73 ) );
  INV_X1 \nop_mux/U71  ( .A(\nop_mux/n67 ), .ZN(\nop_mux/n69 ) );
  AOI22_X1 \nop_mux/U70  ( .A1(operandA_resolved[3]), .A2(\nop_mux/n69 ), .B1(
        1'b0), .B2(\nop_mux/n71 ), .ZN(\nop_mux/n94 ) );
  INV_X1 \nop_mux/U69  ( .A(\nop_mux/n94 ), .ZN(alu_operand[3]) );
  AOI22_X1 \nop_mux/U68  ( .A1(operandA_resolved[26]), .A2(\nop_mux/n68 ), 
        .B1(1'b0), .B2(\nop_mux/n70 ), .ZN(\nop_mux/n88 ) );
  INV_X1 \nop_mux/U67  ( .A(\nop_mux/n88 ), .ZN(alu_operand[26]) );
  AOI22_X1 \nop_mux/U66  ( .A1(operandA_resolved[27]), .A2(\nop_mux/n68 ), 
        .B1(1'b0), .B2(\nop_mux/n70 ), .ZN(\nop_mux/n89 ) );
  INV_X1 \nop_mux/U65  ( .A(\nop_mux/n89 ), .ZN(alu_operand[27]) );
  AOI22_X1 \nop_mux/U64  ( .A1(operandA_resolved[25]), .A2(\nop_mux/n68 ), 
        .B1(1'b0), .B2(\nop_mux/n71 ), .ZN(\nop_mux/n87 ) );
  INV_X1 \nop_mux/U63  ( .A(\nop_mux/n87 ), .ZN(alu_operand[25]) );
  AOI22_X1 \nop_mux/U62  ( .A1(operandA_resolved[24]), .A2(\nop_mux/n68 ), 
        .B1(1'b0), .B2(\nop_mux/n70 ), .ZN(\nop_mux/n86 ) );
  INV_X1 \nop_mux/U61  ( .A(\nop_mux/n86 ), .ZN(alu_operand[24]) );
  AOI22_X1 \nop_mux/U60  ( .A1(operandA_resolved[23]), .A2(\nop_mux/n68 ), 
        .B1(1'b0), .B2(\nop_mux/n71 ), .ZN(\nop_mux/n85 ) );
  INV_X1 \nop_mux/U59  ( .A(\nop_mux/n85 ), .ZN(alu_operand[23]) );
  AOI22_X1 \nop_mux/U58  ( .A1(operandA_resolved[31]), .A2(\nop_mux/n69 ), 
        .B1(1'b0), .B2(\nop_mux/n71 ), .ZN(\nop_mux/n93 ) );
  INV_X1 \nop_mux/U57  ( .A(\nop_mux/n93 ), .ZN(alu_operand[31]) );
  AOI22_X1 \nop_mux/U56  ( .A1(operandA_resolved[19]), .A2(\nop_mux/n68 ), 
        .B1(1'b0), .B2(\nop_mux/n70 ), .ZN(\nop_mux/n81 ) );
  INV_X1 \nop_mux/U55  ( .A(\nop_mux/n81 ), .ZN(alu_operand[19]) );
  AOI22_X1 \nop_mux/U54  ( .A1(operandA_resolved[22]), .A2(\nop_mux/n68 ), 
        .B1(1'b0), .B2(\nop_mux/n70 ), .ZN(\nop_mux/n84 ) );
  INV_X1 \nop_mux/U53  ( .A(\nop_mux/n84 ), .ZN(alu_operand[22]) );
  AOI22_X1 \nop_mux/U52  ( .A1(operandA_resolved[30]), .A2(\nop_mux/n68 ), 
        .B1(1'b0), .B2(\nop_mux/n70 ), .ZN(\nop_mux/n92 ) );
  INV_X1 \nop_mux/U51  ( .A(\nop_mux/n92 ), .ZN(alu_operand[30]) );
  AOI22_X1 \nop_mux/U50  ( .A1(operandA_resolved[16]), .A2(\nop_mux/n68 ), 
        .B1(1'b0), .B2(\nop_mux/n71 ), .ZN(\nop_mux/n78 ) );
  INV_X1 \nop_mux/U49  ( .A(\nop_mux/n78 ), .ZN(alu_operand[16]) );
  AOI22_X1 \nop_mux/U48  ( .A1(operandA_resolved[20]), .A2(\nop_mux/n68 ), 
        .B1(1'b0), .B2(\nop_mux/n70 ), .ZN(\nop_mux/n82 ) );
  INV_X1 \nop_mux/U47  ( .A(\nop_mux/n82 ), .ZN(alu_operand[20]) );
  AOI22_X1 \nop_mux/U46  ( .A1(operandA_resolved[21]), .A2(\nop_mux/n68 ), 
        .B1(1'b0), .B2(\nop_mux/n71 ), .ZN(\nop_mux/n83 ) );
  INV_X1 \nop_mux/U45  ( .A(\nop_mux/n83 ), .ZN(alu_operand[21]) );
  AOI22_X1 \nop_mux/U44  ( .A1(operandA_resolved[28]), .A2(\nop_mux/n68 ), 
        .B1(1'b0), .B2(\nop_mux/n71 ), .ZN(\nop_mux/n90 ) );
  INV_X1 \nop_mux/U43  ( .A(\nop_mux/n90 ), .ZN(alu_operand[28]) );
  AOI22_X1 \nop_mux/U42  ( .A1(operandA_resolved[29]), .A2(\nop_mux/n68 ), 
        .B1(1'b0), .B2(\nop_mux/n70 ), .ZN(\nop_mux/n91 ) );
  INV_X1 \nop_mux/U41  ( .A(\nop_mux/n91 ), .ZN(alu_operand[29]) );
  AOI22_X1 \nop_mux/U40  ( .A1(operandA_resolved[18]), .A2(\nop_mux/n68 ), 
        .B1(1'b0), .B2(\nop_mux/n70 ), .ZN(\nop_mux/n80 ) );
  INV_X1 \nop_mux/U39  ( .A(\nop_mux/n80 ), .ZN(alu_operand[18]) );
  AOI22_X1 \nop_mux/U38  ( .A1(operandA_resolved[17]), .A2(\nop_mux/n68 ), 
        .B1(1'b0), .B2(\nop_mux/n71 ), .ZN(\nop_mux/n79 ) );
  INV_X1 \nop_mux/U37  ( .A(\nop_mux/n79 ), .ZN(alu_operand[17]) );
  AOI22_X1 \nop_mux/U36  ( .A1(operandA_resolved[6]), .A2(\nop_mux/n69 ), .B1(
        1'b0), .B2(\nop_mux/n70 ), .ZN(\nop_mux/n97 ) );
  INV_X1 \nop_mux/U35  ( .A(\nop_mux/n97 ), .ZN(alu_operand[6]) );
  AOI22_X1 \nop_mux/U34  ( .A1(operandA_resolved[9]), .A2(\nop_mux/n69 ), .B1(
        \nop_mux/n71 ), .B2(1'b0), .ZN(\nop_mux/n100 ) );
  INV_X1 \nop_mux/U33  ( .A(\nop_mux/n100 ), .ZN(alu_operand[9]) );
  AOI22_X1 \nop_mux/U32  ( .A1(operandA_resolved[10]), .A2(\nop_mux/n68 ), 
        .B1(1'b0), .B2(\nop_mux/n71 ), .ZN(\nop_mux/n72 ) );
  INV_X1 \nop_mux/U31  ( .A(\nop_mux/n72 ), .ZN(alu_operand[10]) );
  AOI22_X1 \nop_mux/U30  ( .A1(operandA_resolved[12]), .A2(\nop_mux/n68 ), 
        .B1(1'b0), .B2(\nop_mux/n70 ), .ZN(\nop_mux/n74 ) );
  INV_X1 \nop_mux/U29  ( .A(\nop_mux/n74 ), .ZN(alu_operand[12]) );
  AOI22_X1 \nop_mux/U28  ( .A1(operandA_resolved[13]), .A2(\nop_mux/n68 ), 
        .B1(1'b0), .B2(\nop_mux/n70 ), .ZN(\nop_mux/n75 ) );
  INV_X1 \nop_mux/U27  ( .A(\nop_mux/n75 ), .ZN(alu_operand[13]) );
  AOI22_X1 \nop_mux/U26  ( .A1(operandA_resolved[15]), .A2(\nop_mux/n68 ), 
        .B1(1'b0), .B2(\nop_mux/n70 ), .ZN(\nop_mux/n77 ) );
  INV_X1 \nop_mux/U25  ( .A(\nop_mux/n77 ), .ZN(alu_operand[15]) );
  AOI22_X1 \nop_mux/U24  ( .A1(operandA_resolved[4]), .A2(\nop_mux/n69 ), .B1(
        1'b0), .B2(\nop_mux/n71 ), .ZN(\nop_mux/n95 ) );
  INV_X1 \nop_mux/U23  ( .A(\nop_mux/n95 ), .ZN(alu_operand[4]) );
  AOI22_X1 \nop_mux/U22  ( .A1(operandA_resolved[5]), .A2(\nop_mux/n69 ), .B1(
        1'b0), .B2(\nop_mux/n70 ), .ZN(\nop_mux/n96 ) );
  INV_X1 \nop_mux/U21  ( .A(\nop_mux/n96 ), .ZN(alu_operand[5]) );
  AOI22_X1 \nop_mux/U20  ( .A1(operandA_resolved[8]), .A2(\nop_mux/n69 ), .B1(
        1'b0), .B2(\nop_mux/n70 ), .ZN(\nop_mux/n99 ) );
  INV_X1 \nop_mux/U19  ( .A(\nop_mux/n99 ), .ZN(alu_operand[8]) );
  AOI22_X1 \nop_mux/U18  ( .A1(operandA_resolved[7]), .A2(\nop_mux/n69 ), .B1(
        1'b0), .B2(\nop_mux/n70 ), .ZN(\nop_mux/n98 ) );
  INV_X1 \nop_mux/U17  ( .A(\nop_mux/n98 ), .ZN(alu_operand[7]) );
  AOI22_X1 \nop_mux/U16  ( .A1(operandA_resolved[11]), .A2(\nop_mux/n68 ), 
        .B1(1'b0), .B2(\nop_mux/n71 ), .ZN(\nop_mux/n73 ) );
  INV_X1 \nop_mux/U15  ( .A(\nop_mux/n73 ), .ZN(alu_operand[11]) );
  AOI22_X1 \nop_mux/U14  ( .A1(operandA_resolved[14]), .A2(\nop_mux/n68 ), 
        .B1(1'b0), .B2(\nop_mux/n70 ), .ZN(\nop_mux/n76 ) );
  INV_X1 \nop_mux/U13  ( .A(\nop_mux/n76 ), .ZN(alu_operand[14]) );
  INV_X1 \nop_mux/U12  ( .A(\nop_mux/n71 ), .ZN(\nop_mux/n68 ) );
  MUX2_X1 \nop_mux/U11  ( .A(operandA_resolved[1]), .B(1'b0), .S(nop), .Z(
        alu_operand[1]) );
  NAND2_X1 \nop_mux/U10  ( .A1(\nop_mux/n65 ), .A2(\nop_mux/n66 ), .ZN(
        alu_operand[0]) );
  NAND2_X1 \nop_mux/U9  ( .A1(1'b0), .A2(nop), .ZN(\nop_mux/n66 ) );
  NAND2_X1 \nop_mux/U8  ( .A1(operandA_resolved[0]), .A2(\nop_mux/n33 ), .ZN(
        \nop_mux/n65 ) );
  NAND2_X1 \nop_mux/U7  ( .A1(\nop_mux/n43 ), .A2(\nop_mux/n54 ), .ZN(
        alu_operand[2]) );
  NAND2_X1 \nop_mux/U6  ( .A1(1'b0), .A2(nop), .ZN(\nop_mux/n54 ) );
  NAND2_X1 \nop_mux/U5  ( .A1(operandA_resolved[2]), .A2(\nop_mux/n33 ), .ZN(
        \nop_mux/n43 ) );
  INV_X1 \nop_mux/U4  ( .A(nop), .ZN(\nop_mux/n33 ) );
  CLKBUF_X1 \nop_mux/U3  ( .A(nop), .Z(\nop_mux/n67 ) );
  CLKBUF_X2 \nop_mux/U2  ( .A(\nop_mux/n67 ), .Z(\nop_mux/n71 ) );
  BUF_X1 \nop_mux/U1  ( .A(\nop_mux/n67 ), .Z(\nop_mux/n70 ) );
  CLKBUF_X1 \adder/U9  ( .A(\adder/n11 ), .Z(\adder/n18 ) );
  AND2_X1 \adder/U8  ( .A1(\adder/p2 ), .A2(\adder/n13 ), .ZN(\adder/n17 ) );
  AND2_X1 \adder/U7  ( .A1(\adder/p0 ), .A2(n629), .ZN(\adder/n16 ) );
  AND2_X1 \adder/U6  ( .A1(\adder/p1 ), .A2(\adder/n18 ), .ZN(\adder/n15 ) );
  OR2_X1 \adder/U5  ( .A1(\adder/n15 ), .A2(\adder/n10 ), .ZN(\adder/n13 ) );
  OR2_X1 \adder/U4  ( .A1(\adder/g0 ), .A2(\adder/n16 ), .ZN(\adder/n11 ) );
  OR2_X1 \adder/U3  ( .A1(\adder/g2 ), .A2(\adder/n17 ), .ZN(\adder/n14 ) );
  CLKBUF_X1 \adder/U2  ( .A(\adder/g1 ), .Z(\adder/n10 ) );
  OR2_X1 \adder/U1  ( .A1(\adder/g1 ), .A2(\adder/n15 ), .ZN(\adder/n12 ) );
  OAI21_X1 \adder/adder1/U87  ( .B1(\adder/adder1/n50 ), .B2(
        \adder/adder1/n48 ), .A(\adder/adder1/n59 ), .ZN(\adder/adder1/n46 )
         );
  INV_X1 \adder/adder1/U86  ( .A(\adder/adder1/n81 ), .ZN(\adder/adder1/n14 )
         );
  OAI21_X1 \adder/adder1/U85  ( .B1(SYNOPSYS_UNCONNECTED_64), .B2(
        \adder/adder1/n53 ), .A(n629), .ZN(\adder/adder1/n52 ) );
  OAI21_X1 \adder/adder1/U84  ( .B1(SYNOPSYS_UNCONNECTED_57), .B2(
        \adder/adder1/n29 ), .A(\adder/adder1/n82 ), .ZN(\adder/adder1/n28 )
         );
  OAI22_X1 \adder/adder1/U83  ( .A1(\adder/adder1/n14 ), .A2(
        \adder/adder1/n44 ), .B1(\adder/adder1/n45 ), .B2(\adder/adder1/n81 ), 
        .ZN(adder_out[2]) );
  OAI21_X1 \adder/adder1/U82  ( .B1(\adder/adder1/n26 ), .B2(
        \adder/adder1/n82 ), .A(\adder/adder1/n28 ), .ZN(adder_out[7]) );
  XNOR2_X1 \adder/adder1/U81  ( .A(\adder/adder1/n85 ), .B(\adder/adder1/n82 ), 
        .ZN(\adder/adder1/overflow ) );
  AOI21_X1 \adder/adder1/U80  ( .B1(\adder/adder1/n86 ), .B2(n629), .A(
        \adder/adder1/n88 ), .ZN(\adder/adder1/n48 ) );
  NAND4_X1 \adder/adder1/U79  ( .A1(\adder/adder1/n15 ), .A2(
        SYNOPSYS_UNCONNECTED_32), .A3(SYNOPSYS_UNCONNECTED_31), .A4(
        SYNOPSYS_UNCONNECTED_30), .ZN(\adder/adder1/n55 ) );
  OAI21_X1 \adder/adder1/U78  ( .B1(SYNOPSYS_UNCONNECTED_60), .B2(
        \adder/adder1/n40 ), .A(\adder/adder1/n80 ), .ZN(\adder/adder1/n39 )
         );
  OAI21_X1 \adder/adder1/U77  ( .B1(\adder/adder1/n37 ), .B2(
        \adder/adder1/n80 ), .A(\adder/adder1/n39 ), .ZN(adder_out[4]) );
  INV_X1 \adder/adder1/U76  ( .A(\adder/adder1/n34 ), .ZN(\adder/adder1/n13 )
         );
  OAI22_X1 \adder/adder1/U75  ( .A1(\adder/adder1/n33 ), .A2(
        \adder/adder1/n78 ), .B1(\adder/adder1/n77 ), .B2(\adder/adder1/n35 ), 
        .ZN(adder_out[5]) );
  OAI21_X1 \adder/adder1/U74  ( .B1(n629), .B2(\adder/adder1/n51 ), .A(
        \adder/adder1/n52 ), .ZN(adder_out[0]) );
  OAI21_X1 \adder/adder1/U73  ( .B1(\adder/adder1/n30 ), .B2(
        \adder/adder1/n32 ), .A(\adder/adder1/n57 ), .ZN(\adder/adder1/n27 )
         );
  XNOR2_X1 \adder/adder1/U72  ( .A(\adder/adder1/n75 ), .B(\adder/adder1/n31 ), 
        .ZN(adder_out[6]) );
  NOR2_X1 \adder/adder1/U71  ( .A1(\adder/adder1/n87 ), .A2(\adder/adder1/n47 ), .ZN(\adder/adder1/n44 ) );
  AND2_X1 \adder/adder1/U70  ( .A1(alu_operand[2]), .A2(n_2_net__2_), .ZN(
        \adder/adder1/n87 ) );
  XNOR2_X1 \adder/adder1/U69  ( .A(n_2_net__2_), .B(\adder/adder1/n74 ), .ZN(
        \adder/adder1/n45 ) );
  AOI21_X1 \adder/adder1/U68  ( .B1(\adder/adder1/n38 ), .B2(
        SYNOPSYS_UNCONNECTED_28), .A(SYNOPSYS_UNCONNECTED_60), .ZN(
        \adder/adder1/n34 ) );
  OAI21_X1 \adder/adder1/U67  ( .B1(\adder/adder1/n41 ), .B2(
        \adder/adder1/n43 ), .A(\adder/adder1/n58 ), .ZN(\adder/adder1/n38 )
         );
  AND2_X1 \adder/adder1/U66  ( .A1(alu_operand[0]), .A2(n_2_net__0_), .ZN(
        \adder/adder1/n88 ) );
  XNOR2_X1 \adder/adder1/U65  ( .A(n_2_net__0_), .B(\adder/adder1/n79 ), .ZN(
        \adder/adder1/n51 ) );
  OR2_X1 \adder/adder1/U64  ( .A1(alu_operand[0]), .A2(n_2_net__0_), .ZN(
        \adder/adder1/n86 ) );
  NAND2_X1 \adder/adder1/U63  ( .A1(alu_operand[1]), .A2(n_2_net__1_), .ZN(
        \adder/adder1/n59 ) );
  INV_X1 \adder/adder1/U62  ( .A(\adder/adder1/n84 ), .ZN(\adder/adder1/n85 )
         );
  CLKBUF_X1 \adder/adder1/U61  ( .A(\adder/g0 ), .Z(\adder/adder1/n84 ) );
  NOR2_X1 \adder/adder1/U60  ( .A1(alu_operand[1]), .A2(n_2_net__1_), .ZN(
        \adder/adder1/n50 ) );
  AOI21_X1 \adder/adder1/U59  ( .B1(\adder/adder1/n46 ), .B2(
        \adder/adder1/n72 ), .A(\adder/adder1/n87 ), .ZN(\adder/adder1/n41 )
         );
  XNOR2_X1 \adder/adder1/U58  ( .A(\adder/adder1/n71 ), .B(\adder/adder1/n42 ), 
        .ZN(adder_out[3]) );
  XNOR2_X1 \adder/adder1/U57  ( .A(n_2_net__4_), .B(alu_operand[4]), .ZN(
        \adder/adder1/n37 ) );
  XNOR2_X1 \adder/adder1/U56  ( .A(n_2_net__7_), .B(alu_operand[7]), .ZN(
        \adder/adder1/n26 ) );
  NOR2_X1 \adder/adder1/U55  ( .A1(SYNOPSYS_UNCONNECTED_59), .A2(
        \adder/adder1/n36 ), .ZN(\adder/adder1/n35 ) );
  XNOR2_X1 \adder/adder1/U54  ( .A(n_2_net__5_), .B(alu_operand[5]), .ZN(
        \adder/adder1/n33 ) );
  AND2_X1 \adder/adder1/U53  ( .A1(alu_operand[4]), .A2(n_2_net__4_), .ZN(
        SYNOPSYS_UNCONNECTED_60) );
  AND2_X1 \adder/adder1/U52  ( .A1(n_2_net__7_), .A2(alu_operand[7]), .ZN(
        SYNOPSYS_UNCONNECTED_57) );
  AND2_X1 \adder/adder1/U51  ( .A1(alu_operand[5]), .A2(n_2_net__5_), .ZN(
        SYNOPSYS_UNCONNECTED_59) );
  NAND2_X1 \adder/adder1/U50  ( .A1(alu_operand[6]), .A2(n_2_net__6_), .ZN(
        \adder/adder1/n57 ) );
  NAND2_X1 \adder/adder1/U49  ( .A1(alu_operand[3]), .A2(n_2_net__3_), .ZN(
        \adder/adder1/n58 ) );
  NOR2_X1 \adder/adder1/U48  ( .A1(\adder/adder1/n54 ), .A2(\adder/adder1/n55 ), .ZN(\adder/p0 ) );
  NOR2_X1 \adder/adder1/U47  ( .A1(alu_operand[7]), .A2(n_2_net__7_), .ZN(
        \adder/adder1/n29 ) );
  NOR2_X1 \adder/adder1/U46  ( .A1(n_2_net__3_), .A2(alu_operand[3]), .ZN(
        \adder/adder1/n43 ) );
  INV_X1 \adder/adder1/U45  ( .A(\adder/adder1/n57 ), .ZN(
        SYNOPSYS_UNCONNECTED_58) );
  INV_X1 \adder/adder1/U44  ( .A(\adder/adder1/n58 ), .ZN(
        SYNOPSYS_UNCONNECTED_61) );
  INV_X1 \adder/adder1/U43  ( .A(\adder/adder1/n29 ), .ZN(
        SYNOPSYS_UNCONNECTED_25) );
  INV_X1 \adder/adder1/U42  ( .A(\adder/adder1/n36 ), .ZN(
        SYNOPSYS_UNCONNECTED_27) );
  INV_X1 \adder/adder1/U41  ( .A(\adder/adder1/n32 ), .ZN(
        SYNOPSYS_UNCONNECTED_26) );
  NOR2_X1 \adder/adder1/U40  ( .A1(SYNOPSYS_UNCONNECTED_61), .A2(
        \adder/adder1/n70 ), .ZN(\adder/adder1/n42 ) );
  OR2_X1 \adder/adder1/U39  ( .A1(SYNOPSYS_UNCONNECTED_63), .A2(
        \adder/adder1/n69 ), .ZN(\adder/adder1/n83 ) );
  XOR2_X1 \adder/adder1/U38  ( .A(\adder/adder1/n68 ), .B(\adder/adder1/n83 ), 
        .Z(adder_out[1]) );
  NOR2_X1 \adder/adder1/U37  ( .A1(SYNOPSYS_UNCONNECTED_58), .A2(
        \adder/adder1/n32 ), .ZN(\adder/adder1/n31 ) );
  INV_X1 \adder/adder1/U36  ( .A(SYNOPSYS_UNCONNECTED_32), .ZN(
        \adder/adder1/n53 ) );
  INV_X1 \adder/adder1/U35  ( .A(\adder/adder1/n29 ), .ZN(\adder/adder1/n15 )
         );
  INV_X1 \adder/adder1/U34  ( .A(\adder/adder1/n32 ), .ZN(\adder/adder1/n17 )
         );
  NAND4_X1 \adder/adder1/U33  ( .A1(SYNOPSYS_UNCONNECTED_29), .A2(
        SYNOPSYS_UNCONNECTED_28), .A3(\adder/adder1/n62 ), .A4(
        \adder/adder1/n17 ), .ZN(\adder/adder1/n54 ) );
  AOI21_X1 \adder/adder1/U32  ( .B1(\adder/adder1/n13 ), .B2(
        \adder/adder1/n62 ), .A(SYNOPSYS_UNCONNECTED_59), .ZN(
        \adder/adder1/n30 ) );
  CLKBUF_X1 \adder/adder1/U31  ( .A(\adder/adder1/n27 ), .Z(\adder/adder1/n82 ) );
  CLKBUF_X1 \adder/adder1/U30  ( .A(\adder/adder1/n46 ), .Z(\adder/adder1/n81 ) );
  CLKBUF_X1 \adder/adder1/U29  ( .A(\adder/adder1/n38 ), .Z(\adder/adder1/n80 ) );
  CLKBUF_X1 \adder/adder1/U28  ( .A(alu_operand[0]), .Z(\adder/adder1/n79 ) );
  CLKBUF_X1 \adder/adder1/U27  ( .A(\adder/adder1/n13 ), .Z(\adder/adder1/n78 ) );
  INV_X1 \adder/adder1/U26  ( .A(\adder/adder1/n78 ), .ZN(\adder/adder1/n77 )
         );
  OR2_X1 \adder/adder1/U25  ( .A1(\adder/adder1/n60 ), .A2(n_2_net__1_), .ZN(
        SYNOPSYS_UNCONNECTED_31) );
  AOI21_X1 \adder/adder1/U24  ( .B1(\adder/adder1/n78 ), .B2(
        SYNOPSYS_UNCONNECTED_27), .A(SYNOPSYS_UNCONNECTED_59), .ZN(
        \adder/adder1/n75 ) );
  CLKBUF_X1 \adder/adder1/U23  ( .A(alu_operand[2]), .Z(\adder/adder1/n74 ) );
  OR2_X1 \adder/adder1/U22  ( .A1(alu_operand[4]), .A2(n_2_net__4_), .ZN(
        SYNOPSYS_UNCONNECTED_28) );
  INV_X1 \adder/adder1/U21  ( .A(SYNOPSYS_UNCONNECTED_28), .ZN(
        \adder/adder1/n40 ) );
  OR2_X1 \adder/adder1/U20  ( .A1(alu_operand[2]), .A2(n_2_net__2_), .ZN(
        \adder/adder1/n72 ) );
  INV_X1 \adder/adder1/U19  ( .A(SYNOPSYS_UNCONNECTED_30), .ZN(
        \adder/adder1/n47 ) );
  AOI21_X1 \adder/adder1/U18  ( .B1(\adder/adder1/n81 ), .B2(
        SYNOPSYS_UNCONNECTED_30), .A(\adder/adder1/n87 ), .ZN(
        \adder/adder1/n71 ) );
  INV_X1 \adder/adder1/U17  ( .A(SYNOPSYS_UNCONNECTED_29), .ZN(
        \adder/adder1/n70 ) );
  INV_X1 \adder/adder1/U16  ( .A(\adder/adder1/n49 ), .ZN(
        SYNOPSYS_UNCONNECTED_63) );
  INV_X1 \adder/adder1/U15  ( .A(SYNOPSYS_UNCONNECTED_31), .ZN(
        \adder/adder1/n69 ) );
  AOI21_X1 \adder/adder1/U14  ( .B1(SYNOPSYS_UNCONNECTED_32), .B2(n629), .A(
        SYNOPSYS_UNCONNECTED_64), .ZN(\adder/adder1/n68 ) );
  OR2_X1 \adder/adder1/U13  ( .A1(alu_operand[3]), .A2(n_2_net__3_), .ZN(
        SYNOPSYS_UNCONNECTED_29) );
  CLKBUF_X1 \adder/adder1/U12  ( .A(\adder/adder1/n87 ), .Z(
        SYNOPSYS_UNCONNECTED_62) );
  CLKBUF_X1 \adder/adder1/U11  ( .A(\adder/adder1/n88 ), .Z(
        SYNOPSYS_UNCONNECTED_64) );
  INV_X1 \adder/adder1/U10  ( .A(SYNOPSYS_UNCONNECTED_57), .ZN(
        \adder/adder1/n64 ) );
  INV_X1 \adder/adder1/U9  ( .A(\adder/adder1/n27 ), .ZN(\adder/adder1/n63 )
         );
  OAI21_X1 \adder/adder1/U8  ( .B1(\adder/adder1/n63 ), .B2(\adder/adder1/n29 ), .A(\adder/adder1/n64 ), .ZN(\adder/g0 ) );
  OR2_X1 \adder/adder1/U7  ( .A1(alu_operand[5]), .A2(n_2_net__5_), .ZN(
        \adder/adder1/n62 ) );
  CLKBUF_X1 \adder/adder1/U6  ( .A(\adder/adder1/n72 ), .Z(
        SYNOPSYS_UNCONNECTED_30) );
  NOR2_X1 \adder/adder1/U5  ( .A1(alu_operand[6]), .A2(n_2_net__6_), .ZN(
        \adder/adder1/n32 ) );
  CLKBUF_X1 \adder/adder1/U4  ( .A(alu_operand[1]), .Z(\adder/adder1/n60 ) );
  INV_X1 \adder/adder1/U3  ( .A(\adder/adder1/n62 ), .ZN(\adder/adder1/n36 )
         );
  OR2_X1 \adder/adder1/U2  ( .A1(alu_operand[0]), .A2(n_2_net__0_), .ZN(
        SYNOPSYS_UNCONNECTED_32) );
  CLKBUF_X1 \adder/adder1/U1  ( .A(\adder/adder1/n59 ), .Z(\adder/adder1/n49 )
         );
  OAI21_X1 \adder/adder2/U78  ( .B1(SYNOPSYS_UNCONNECTED_49), .B2(
        \adder/adder2/n104 ), .A(\adder/adder2/n106 ), .ZN(\adder/adder2/n105 ) );
  OAI21_X1 \adder/adder2/U77  ( .B1(SYNOPSYS_UNCONNECTED_52), .B2(
        \adder/adder2/n93 ), .A(\adder/adder2/n72 ), .ZN(\adder/adder2/n94 )
         );
  INV_X1 \adder/adder2/U76  ( .A(\adder/adder2/n73 ), .ZN(\adder/adder2/n109 )
         );
  OAI22_X1 \adder/adder2/U75  ( .A1(\adder/adder2/n109 ), .A2(
        \adder/adder2/n89 ), .B1(\adder/adder2/n88 ), .B2(\adder/adder2/n73 ), 
        .ZN(adder_out[10]) );
  OAI21_X1 \adder/adder2/U74  ( .B1(\adder/adder2/n107 ), .B2(
        \adder/adder2/n106 ), .A(\adder/adder2/n105 ), .ZN(adder_out[15]) );
  OAI21_X1 \adder/adder2/U73  ( .B1(\adder/adder2/n96 ), .B2(
        \adder/adder2/n72 ), .A(\adder/adder2/n94 ), .ZN(adder_out[12]) );
  XNOR2_X1 \adder/adder2/U72  ( .A(\adder/adder2/n74 ), .B(\adder/adder2/n106 ), .ZN(\adder/adder2/overflow ) );
  OAI21_X1 \adder/adder2/U71  ( .B1(\adder/adder2/n85 ), .B2(
        \adder/adder2/n83 ), .A(\adder/adder2/n75 ), .ZN(\adder/adder2/n87 )
         );
  OAI21_X1 \adder/adder2/U70  ( .B1(\adder/adder2/n103 ), .B2(
        \adder/adder2/n101 ), .A(\adder/adder2/n77 ), .ZN(\adder/adder2/n106 )
         );
  XNOR2_X1 \adder/adder2/U69  ( .A(\adder/adder2/n68 ), .B(\adder/adder2/n84 ), 
        .ZN(adder_out[9]) );
  XNOR2_X1 \adder/adder2/U68  ( .A(\adder/adder2/n71 ), .B(\adder/adder2/n102 ), .ZN(adder_out[14]) );
  AOI21_X1 \adder/adder2/U67  ( .B1(\adder/n11 ), .B2(SYNOPSYS_UNCONNECTED_24), 
        .A(SYNOPSYS_UNCONNECTED_56), .ZN(\adder/adder2/n85 ) );
  OAI21_X1 \adder/adder2/U66  ( .B1(\adder/adder2/n92 ), .B2(
        \adder/adder2/n90 ), .A(\adder/adder2/n76 ), .ZN(\adder/adder2/n95 )
         );
  XNOR2_X1 \adder/adder2/U65  ( .A(\adder/adder2/n69 ), .B(\adder/adder2/n91 ), 
        .ZN(adder_out[11]) );
  AOI21_X1 \adder/adder2/U64  ( .B1(\adder/adder2/n87 ), .B2(
        SYNOPSYS_UNCONNECTED_22), .A(SYNOPSYS_UNCONNECTED_54), .ZN(
        \adder/adder2/n92 ) );
  AOI21_X1 \adder/adder2/U63  ( .B1(\adder/adder2/n95 ), .B2(
        SYNOPSYS_UNCONNECTED_20), .A(SYNOPSYS_UNCONNECTED_52), .ZN(
        \adder/adder2/n99 ) );
  INV_X1 \adder/adder2/U62  ( .A(\adder/adder2/n67 ), .ZN(\adder/adder2/n110 )
         );
  OAI22_X1 \adder/adder2/U61  ( .A1(\adder/adder2/n100 ), .A2(
        \adder/adder2/n110 ), .B1(\adder/adder2/n70 ), .B2(\adder/adder2/n98 ), 
        .ZN(adder_out[13]) );
  OAI21_X1 \adder/adder2/U60  ( .B1(SYNOPSYS_UNCONNECTED_56), .B2(
        \adder/adder2/n80 ), .A(\adder/adder2/n65 ), .ZN(\adder/adder2/n81 )
         );
  OAI21_X1 \adder/adder2/U59  ( .B1(\adder/adder2/n65 ), .B2(
        \adder/adder2/n82 ), .A(\adder/adder2/n81 ), .ZN(adder_out[8]) );
  INV_X1 \adder/adder2/U58  ( .A(\adder/adder2/n66 ), .ZN(\adder/adder2/n74 )
         );
  AND2_X1 \adder/adder2/U57  ( .A1(n_2_net__15_), .A2(alu_operand[15]), .ZN(
        SYNOPSYS_UNCONNECTED_49) );
  NAND2_X1 \adder/adder2/U56  ( .A1(alu_operand[14]), .A2(n_2_net__14_), .ZN(
        \adder/adder2/n77 ) );
  XNOR2_X1 \adder/adder2/U55  ( .A(n_2_net__8_), .B(alu_operand[8]), .ZN(
        \adder/adder2/n82 ) );
  XNOR2_X1 \adder/adder2/U54  ( .A(n_2_net__15_), .B(alu_operand[15]), .ZN(
        \adder/adder2/n107 ) );
  XNOR2_X1 \adder/adder2/U53  ( .A(n_2_net__12_), .B(alu_operand[12]), .ZN(
        \adder/adder2/n96 ) );
  NOR2_X1 \adder/adder2/U52  ( .A1(SYNOPSYS_UNCONNECTED_54), .A2(
        \adder/adder2/n86 ), .ZN(\adder/adder2/n89 ) );
  XNOR2_X1 \adder/adder2/U51  ( .A(n_2_net__10_), .B(alu_operand[10]), .ZN(
        \adder/adder2/n88 ) );
  NOR2_X1 \adder/adder2/U50  ( .A1(SYNOPSYS_UNCONNECTED_51), .A2(
        \adder/adder2/n97 ), .ZN(\adder/adder2/n98 ) );
  XNOR2_X1 \adder/adder2/U49  ( .A(n_2_net__13_), .B(alu_operand[13]), .ZN(
        \adder/adder2/n100 ) );
  AND2_X1 \adder/adder2/U48  ( .A1(alu_operand[12]), .A2(n_2_net__12_), .ZN(
        SYNOPSYS_UNCONNECTED_52) );
  AND2_X1 \adder/adder2/U47  ( .A1(alu_operand[8]), .A2(n_2_net__8_), .ZN(
        SYNOPSYS_UNCONNECTED_56) );
  AND2_X1 \adder/adder2/U46  ( .A1(alu_operand[10]), .A2(n_2_net__10_), .ZN(
        SYNOPSYS_UNCONNECTED_54) );
  AND2_X1 \adder/adder2/U45  ( .A1(alu_operand[13]), .A2(n_2_net__13_), .ZN(
        SYNOPSYS_UNCONNECTED_51) );
  NAND2_X1 \adder/adder2/U44  ( .A1(alu_operand[11]), .A2(n_2_net__11_), .ZN(
        \adder/adder2/n76 ) );
  NAND2_X1 \adder/adder2/U43  ( .A1(alu_operand[9]), .A2(n_2_net__9_), .ZN(
        \adder/adder2/n75 ) );
  NOR2_X1 \adder/adder2/U42  ( .A1(alu_operand[12]), .A2(n_2_net__12_), .ZN(
        \adder/adder2/n93 ) );
  NOR2_X1 \adder/adder2/U41  ( .A1(alu_operand[15]), .A2(n_2_net__15_), .ZN(
        \adder/adder2/n104 ) );
  NOR2_X1 \adder/adder2/U40  ( .A1(alu_operand[8]), .A2(n_2_net__8_), .ZN(
        \adder/adder2/n80 ) );
  NOR2_X1 \adder/adder2/U39  ( .A1(alu_operand[10]), .A2(n_2_net__10_), .ZN(
        \adder/adder2/n86 ) );
  NOR2_X1 \adder/adder2/U38  ( .A1(alu_operand[13]), .A2(n_2_net__13_), .ZN(
        \adder/adder2/n97 ) );
  NOR2_X1 \adder/adder2/U37  ( .A1(alu_operand[11]), .A2(n_2_net__11_), .ZN(
        \adder/adder2/n90 ) );
  NOR2_X1 \adder/adder2/U36  ( .A1(alu_operand[14]), .A2(n_2_net__14_), .ZN(
        \adder/adder2/n101 ) );
  NOR2_X1 \adder/adder2/U35  ( .A1(alu_operand[9]), .A2(n_2_net__9_), .ZN(
        \adder/adder2/n83 ) );
  INV_X1 \adder/adder2/U34  ( .A(\adder/adder2/n77 ), .ZN(
        SYNOPSYS_UNCONNECTED_50) );
  INV_X1 \adder/adder2/U33  ( .A(\adder/adder2/n76 ), .ZN(
        SYNOPSYS_UNCONNECTED_53) );
  INV_X1 \adder/adder2/U32  ( .A(\adder/adder2/n75 ), .ZN(
        SYNOPSYS_UNCONNECTED_55) );
  INV_X1 \adder/adder2/U31  ( .A(\adder/adder2/n93 ), .ZN(
        SYNOPSYS_UNCONNECTED_20) );
  INV_X1 \adder/adder2/U30  ( .A(\adder/adder2/n80 ), .ZN(
        SYNOPSYS_UNCONNECTED_24) );
  INV_X1 \adder/adder2/U29  ( .A(\adder/adder2/n97 ), .ZN(
        SYNOPSYS_UNCONNECTED_19) );
  INV_X1 \adder/adder2/U28  ( .A(\adder/adder2/n86 ), .ZN(
        SYNOPSYS_UNCONNECTED_22) );
  INV_X1 \adder/adder2/U27  ( .A(\adder/adder2/n83 ), .ZN(
        SYNOPSYS_UNCONNECTED_23) );
  INV_X1 \adder/adder2/U26  ( .A(\adder/adder2/n101 ), .ZN(
        SYNOPSYS_UNCONNECTED_18) );
  INV_X1 \adder/adder2/U25  ( .A(\adder/adder2/n90 ), .ZN(
        SYNOPSYS_UNCONNECTED_21) );
  NOR2_X1 \adder/adder2/U24  ( .A1(SYNOPSYS_UNCONNECTED_55), .A2(
        \adder/adder2/n83 ), .ZN(\adder/adder2/n84 ) );
  NOR2_X1 \adder/adder2/U23  ( .A1(SYNOPSYS_UNCONNECTED_53), .A2(
        \adder/adder2/n90 ), .ZN(\adder/adder2/n91 ) );
  NOR2_X1 \adder/adder2/U22  ( .A1(SYNOPSYS_UNCONNECTED_50), .A2(
        \adder/adder2/n101 ), .ZN(\adder/adder2/n102 ) );
  INV_X1 \adder/adder2/U21  ( .A(\adder/adder2/n104 ), .ZN(
        SYNOPSYS_UNCONNECTED_17) );
  NAND4_X1 \adder/adder2/U20  ( .A1(SYNOPSYS_UNCONNECTED_21), .A2(
        SYNOPSYS_UNCONNECTED_20), .A3(SYNOPSYS_UNCONNECTED_19), .A4(
        \adder/adder2/n60 ), .ZN(\adder/adder2/n79 ) );
  NAND4_X1 \adder/adder2/U19  ( .A1(SYNOPSYS_UNCONNECTED_17), .A2(
        SYNOPSYS_UNCONNECTED_24), .A3(SYNOPSYS_UNCONNECTED_23), .A4(
        SYNOPSYS_UNCONNECTED_22), .ZN(\adder/adder2/n78 ) );
  NOR2_X1 \adder/adder2/U18  ( .A1(\adder/adder2/n79 ), .A2(\adder/adder2/n78 ), .ZN(\adder/p1 ) );
  CLKBUF_X1 \adder/adder2/U17  ( .A(\adder/adder2/n87 ), .Z(\adder/adder2/n73 ) );
  CLKBUF_X1 \adder/adder2/U16  ( .A(\adder/adder2/n95 ), .Z(\adder/adder2/n72 ) );
  AOI21_X1 \adder/adder2/U15  ( .B1(\adder/adder2/n110 ), .B2(
        SYNOPSYS_UNCONNECTED_19), .A(SYNOPSYS_UNCONNECTED_51), .ZN(
        \adder/adder2/n71 ) );
  INV_X1 \adder/adder2/U14  ( .A(\adder/adder2/n110 ), .ZN(\adder/adder2/n70 )
         );
  AOI21_X1 \adder/adder2/U13  ( .B1(\adder/adder2/n73 ), .B2(
        SYNOPSYS_UNCONNECTED_22), .A(SYNOPSYS_UNCONNECTED_54), .ZN(
        \adder/adder2/n69 ) );
  AOI21_X1 \adder/adder2/U12  ( .B1(\adder/adder2/n65 ), .B2(
        SYNOPSYS_UNCONNECTED_24), .A(SYNOPSYS_UNCONNECTED_56), .ZN(
        \adder/adder2/n68 ) );
  AOI21_X1 \adder/adder2/U11  ( .B1(\adder/adder2/n72 ), .B2(
        SYNOPSYS_UNCONNECTED_20), .A(SYNOPSYS_UNCONNECTED_52), .ZN(
        \adder/adder2/n67 ) );
  CLKBUF_X1 \adder/adder2/U10  ( .A(\adder/g1 ), .Z(\adder/adder2/n66 ) );
  CLKBUF_X1 \adder/adder2/U9  ( .A(\adder/n11 ), .Z(\adder/adder2/n65 ) );
  INV_X1 \adder/adder2/U8  ( .A(\adder/adder2/n56 ), .ZN(\adder/adder2/n103 )
         );
  INV_X1 \adder/adder2/U7  ( .A(SYNOPSYS_UNCONNECTED_51), .ZN(
        \adder/adder2/n63 ) );
  OAI21_X1 \adder/adder2/U6  ( .B1(\adder/adder2/n99 ), .B2(\adder/adder2/n97 ), .A(\adder/adder2/n63 ), .ZN(\adder/adder2/n64 ) );
  INV_X1 \adder/adder2/U5  ( .A(SYNOPSYS_UNCONNECTED_49), .ZN(
        \adder/adder2/n62 ) );
  OAI21_X1 \adder/adder2/U4  ( .B1(\adder/adder2/n61 ), .B2(
        \adder/adder2/n104 ), .A(\adder/adder2/n62 ), .ZN(\adder/g1 ) );
  INV_X1 \adder/adder2/U3  ( .A(\adder/adder2/n101 ), .ZN(\adder/adder2/n60 )
         );
  AOI21_X1 \adder/adder2/U2  ( .B1(\adder/adder2/n64 ), .B2(\adder/adder2/n60 ), .A(SYNOPSYS_UNCONNECTED_50), .ZN(\adder/adder2/n61 ) );
  CLKBUF_X1 \adder/adder2/U1  ( .A(\adder/adder2/n64 ), .Z(\adder/adder2/n56 )
         );
  OAI21_X1 \adder/adder3/U78  ( .B1(SYNOPSYS_UNCONNECTED_41), .B2(
        \adder/adder3/n104 ), .A(\adder/adder3/n106 ), .ZN(\adder/adder3/n105 ) );
  OAI21_X1 \adder/adder3/U77  ( .B1(SYNOPSYS_UNCONNECTED_44), .B2(
        \adder/adder3/n93 ), .A(\adder/adder3/n73 ), .ZN(\adder/adder3/n94 )
         );
  INV_X1 \adder/adder3/U76  ( .A(\adder/adder3/n74 ), .ZN(\adder/adder3/n109 )
         );
  OAI22_X1 \adder/adder3/U75  ( .A1(\adder/adder3/n109 ), .A2(
        \adder/adder3/n89 ), .B1(\adder/adder3/n88 ), .B2(\adder/adder3/n74 ), 
        .ZN(adder_out[18]) );
  OAI21_X1 \adder/adder3/U74  ( .B1(\adder/adder3/n107 ), .B2(
        \adder/adder3/n106 ), .A(\adder/adder3/n105 ), .ZN(adder_out[23]) );
  OAI21_X1 \adder/adder3/U73  ( .B1(\adder/adder3/n96 ), .B2(
        \adder/adder3/n73 ), .A(\adder/adder3/n94 ), .ZN(adder_out[20]) );
  XNOR2_X1 \adder/adder3/U72  ( .A(\adder/adder3/n72 ), .B(\adder/adder3/n106 ), .ZN(\adder/adder3/overflow ) );
  OAI21_X1 \adder/adder3/U71  ( .B1(\adder/adder3/n85 ), .B2(
        \adder/adder3/n83 ), .A(\adder/adder3/n75 ), .ZN(\adder/adder3/n87 )
         );
  XNOR2_X1 \adder/adder3/U70  ( .A(\adder/adder3/n68 ), .B(\adder/adder3/n84 ), 
        .ZN(adder_out[17]) );
  XNOR2_X1 \adder/adder3/U69  ( .A(\adder/adder3/n71 ), .B(\adder/adder3/n102 ), .ZN(adder_out[22]) );
  AOI21_X1 \adder/adder3/U68  ( .B1(\adder/n12 ), .B2(SYNOPSYS_UNCONNECTED_16), 
        .A(SYNOPSYS_UNCONNECTED_48), .ZN(\adder/adder3/n85 ) );
  OAI21_X1 \adder/adder3/U67  ( .B1(\adder/adder3/n92 ), .B2(
        \adder/adder3/n90 ), .A(\adder/adder3/n76 ), .ZN(\adder/adder3/n95 )
         );
  XNOR2_X1 \adder/adder3/U66  ( .A(\adder/adder3/n70 ), .B(\adder/adder3/n91 ), 
        .ZN(adder_out[19]) );
  AOI21_X1 \adder/adder3/U65  ( .B1(\adder/adder3/n87 ), .B2(
        SYNOPSYS_UNCONNECTED_14), .A(SYNOPSYS_UNCONNECTED_46), .ZN(
        \adder/adder3/n92 ) );
  AOI21_X1 \adder/adder3/U64  ( .B1(\adder/adder3/n95 ), .B2(
        SYNOPSYS_UNCONNECTED_12), .A(SYNOPSYS_UNCONNECTED_44), .ZN(
        \adder/adder3/n99 ) );
  INV_X1 \adder/adder3/U63  ( .A(\adder/adder3/n66 ), .ZN(\adder/adder3/n110 )
         );
  OAI22_X1 \adder/adder3/U62  ( .A1(\adder/adder3/n100 ), .A2(
        \adder/adder3/n110 ), .B1(\adder/adder3/n69 ), .B2(\adder/adder3/n98 ), 
        .ZN(adder_out[21]) );
  OAI21_X1 \adder/adder3/U61  ( .B1(SYNOPSYS_UNCONNECTED_48), .B2(
        \adder/adder3/n80 ), .A(\adder/adder3/n65 ), .ZN(\adder/adder3/n81 )
         );
  OAI21_X1 \adder/adder3/U60  ( .B1(\adder/adder3/n82 ), .B2(
        \adder/adder3/n65 ), .A(\adder/adder3/n81 ), .ZN(adder_out[16]) );
  AND2_X1 \adder/adder3/U59  ( .A1(alu_operand[20]), .A2(n_2_net__20_), .ZN(
        SYNOPSYS_UNCONNECTED_44) );
  AND2_X1 \adder/adder3/U58  ( .A1(alu_operand[16]), .A2(n_2_net__16_), .ZN(
        SYNOPSYS_UNCONNECTED_48) );
  AND2_X1 \adder/adder3/U57  ( .A1(n_2_net__23_), .A2(alu_operand[23]), .ZN(
        SYNOPSYS_UNCONNECTED_41) );
  AND2_X1 \adder/adder3/U56  ( .A1(alu_operand[18]), .A2(n_2_net__18_), .ZN(
        SYNOPSYS_UNCONNECTED_46) );
  AND2_X1 \adder/adder3/U55  ( .A1(alu_operand[21]), .A2(n_2_net__21_), .ZN(
        SYNOPSYS_UNCONNECTED_43) );
  NAND2_X1 \adder/adder3/U54  ( .A1(alu_operand[17]), .A2(n_2_net__17_), .ZN(
        \adder/adder3/n75 ) );
  NAND2_X1 \adder/adder3/U53  ( .A1(alu_operand[19]), .A2(n_2_net__19_), .ZN(
        \adder/adder3/n76 ) );
  NAND2_X1 \adder/adder3/U52  ( .A1(alu_operand[22]), .A2(n_2_net__22_), .ZN(
        \adder/adder3/n77 ) );
  NOR2_X1 \adder/adder3/U51  ( .A1(alu_operand[23]), .A2(n_2_net__23_), .ZN(
        \adder/adder3/n104 ) );
  NOR2_X1 \adder/adder3/U50  ( .A1(alu_operand[20]), .A2(n_2_net__20_), .ZN(
        \adder/adder3/n93 ) );
  NOR2_X1 \adder/adder3/U49  ( .A1(alu_operand[16]), .A2(n_2_net__16_), .ZN(
        \adder/adder3/n80 ) );
  NOR2_X1 \adder/adder3/U48  ( .A1(alu_operand[18]), .A2(n_2_net__18_), .ZN(
        \adder/adder3/n86 ) );
  NOR2_X1 \adder/adder3/U47  ( .A1(alu_operand[21]), .A2(n_2_net__21_), .ZN(
        \adder/adder3/n97 ) );
  NOR2_X1 \adder/adder3/U46  ( .A1(alu_operand[19]), .A2(n_2_net__19_), .ZN(
        \adder/adder3/n90 ) );
  NOR2_X1 \adder/adder3/U45  ( .A1(alu_operand[22]), .A2(n_2_net__22_), .ZN(
        \adder/adder3/n101 ) );
  XNOR2_X1 \adder/adder3/U44  ( .A(n_2_net__16_), .B(alu_operand[16]), .ZN(
        \adder/adder3/n82 ) );
  XNOR2_X1 \adder/adder3/U43  ( .A(n_2_net__20_), .B(alu_operand[20]), .ZN(
        \adder/adder3/n96 ) );
  NOR2_X1 \adder/adder3/U42  ( .A1(SYNOPSYS_UNCONNECTED_46), .A2(
        \adder/adder3/n86 ), .ZN(\adder/adder3/n89 ) );
  XNOR2_X1 \adder/adder3/U41  ( .A(n_2_net__18_), .B(alu_operand[18]), .ZN(
        \adder/adder3/n88 ) );
  XNOR2_X1 \adder/adder3/U40  ( .A(n_2_net__23_), .B(alu_operand[23]), .ZN(
        \adder/adder3/n107 ) );
  NOR2_X1 \adder/adder3/U39  ( .A1(SYNOPSYS_UNCONNECTED_43), .A2(
        \adder/adder3/n97 ), .ZN(\adder/adder3/n98 ) );
  XNOR2_X1 \adder/adder3/U38  ( .A(n_2_net__21_), .B(alu_operand[21]), .ZN(
        \adder/adder3/n100 ) );
  INV_X1 \adder/adder3/U37  ( .A(\adder/adder3/n77 ), .ZN(
        SYNOPSYS_UNCONNECTED_42) );
  INV_X1 \adder/adder3/U36  ( .A(\adder/adder3/n76 ), .ZN(
        SYNOPSYS_UNCONNECTED_45) );
  INV_X1 \adder/adder3/U35  ( .A(\adder/adder3/n75 ), .ZN(
        SYNOPSYS_UNCONNECTED_47) );
  INV_X1 \adder/adder3/U34  ( .A(\adder/adder3/n104 ), .ZN(
        SYNOPSYS_UNCONNECTED_9) );
  INV_X1 \adder/adder3/U33  ( .A(\adder/adder3/n93 ), .ZN(
        SYNOPSYS_UNCONNECTED_12) );
  INV_X1 \adder/adder3/U32  ( .A(\adder/adder3/n97 ), .ZN(
        SYNOPSYS_UNCONNECTED_11) );
  INV_X1 \adder/adder3/U31  ( .A(\adder/adder3/n86 ), .ZN(
        SYNOPSYS_UNCONNECTED_14) );
  INV_X1 \adder/adder3/U30  ( .A(\adder/adder3/n83 ), .ZN(
        SYNOPSYS_UNCONNECTED_15) );
  INV_X1 \adder/adder3/U29  ( .A(\adder/adder3/n101 ), .ZN(
        SYNOPSYS_UNCONNECTED_10) );
  INV_X1 \adder/adder3/U28  ( .A(\adder/adder3/n90 ), .ZN(
        SYNOPSYS_UNCONNECTED_13) );
  INV_X1 \adder/adder3/U27  ( .A(\adder/adder3/n80 ), .ZN(
        SYNOPSYS_UNCONNECTED_16) );
  NAND4_X1 \adder/adder3/U26  ( .A1(SYNOPSYS_UNCONNECTED_13), .A2(
        SYNOPSYS_UNCONNECTED_12), .A3(SYNOPSYS_UNCONNECTED_11), .A4(
        \adder/adder3/n60 ), .ZN(\adder/adder3/n79 ) );
  NAND4_X1 \adder/adder3/U25  ( .A1(SYNOPSYS_UNCONNECTED_9), .A2(
        SYNOPSYS_UNCONNECTED_16), .A3(SYNOPSYS_UNCONNECTED_15), .A4(
        SYNOPSYS_UNCONNECTED_14), .ZN(\adder/adder3/n78 ) );
  NOR2_X1 \adder/adder3/U24  ( .A1(SYNOPSYS_UNCONNECTED_47), .A2(
        \adder/adder3/n83 ), .ZN(\adder/adder3/n84 ) );
  NOR2_X1 \adder/adder3/U23  ( .A1(SYNOPSYS_UNCONNECTED_45), .A2(
        \adder/adder3/n90 ), .ZN(\adder/adder3/n91 ) );
  NOR2_X1 \adder/adder3/U22  ( .A1(SYNOPSYS_UNCONNECTED_42), .A2(
        \adder/adder3/n101 ), .ZN(\adder/adder3/n102 ) );
  NOR2_X1 \adder/adder3/U21  ( .A1(\adder/adder3/n79 ), .A2(\adder/adder3/n78 ), .ZN(\adder/p2 ) );
  CLKBUF_X1 \adder/adder3/U20  ( .A(\adder/adder3/n87 ), .Z(\adder/adder3/n74 ) );
  CLKBUF_X1 \adder/adder3/U19  ( .A(\adder/adder3/n95 ), .Z(\adder/adder3/n73 ) );
  INV_X1 \adder/adder3/U18  ( .A(\adder/adder3/n67 ), .ZN(\adder/adder3/n72 )
         );
  AOI21_X1 \adder/adder3/U17  ( .B1(\adder/adder3/n110 ), .B2(
        SYNOPSYS_UNCONNECTED_11), .A(SYNOPSYS_UNCONNECTED_43), .ZN(
        \adder/adder3/n71 ) );
  AOI21_X1 \adder/adder3/U16  ( .B1(\adder/adder3/n74 ), .B2(
        SYNOPSYS_UNCONNECTED_14), .A(SYNOPSYS_UNCONNECTED_46), .ZN(
        \adder/adder3/n70 ) );
  INV_X1 \adder/adder3/U15  ( .A(\adder/adder3/n110 ), .ZN(\adder/adder3/n69 )
         );
  AOI21_X1 \adder/adder3/U14  ( .B1(\adder/adder3/n65 ), .B2(
        SYNOPSYS_UNCONNECTED_16), .A(SYNOPSYS_UNCONNECTED_48), .ZN(
        \adder/adder3/n68 ) );
  CLKBUF_X1 \adder/adder3/U13  ( .A(\adder/g2 ), .Z(\adder/adder3/n67 ) );
  AOI21_X1 \adder/adder3/U12  ( .B1(\adder/adder3/n73 ), .B2(
        SYNOPSYS_UNCONNECTED_12), .A(SYNOPSYS_UNCONNECTED_44), .ZN(
        \adder/adder3/n66 ) );
  CLKBUF_X1 \adder/adder3/U11  ( .A(\adder/n12 ), .Z(\adder/adder3/n65 ) );
  INV_X1 \adder/adder3/U10  ( .A(\adder/adder3/n56 ), .ZN(\adder/adder3/n103 )
         );
  INV_X1 \adder/adder3/U9  ( .A(SYNOPSYS_UNCONNECTED_43), .ZN(
        \adder/adder3/n63 ) );
  OAI21_X1 \adder/adder3/U8  ( .B1(\adder/adder3/n99 ), .B2(\adder/adder3/n97 ), .A(\adder/adder3/n63 ), .ZN(\adder/adder3/n64 ) );
  INV_X1 \adder/adder3/U7  ( .A(SYNOPSYS_UNCONNECTED_41), .ZN(
        \adder/adder3/n62 ) );
  OAI21_X1 \adder/adder3/U6  ( .B1(\adder/adder3/n61 ), .B2(
        \adder/adder3/n104 ), .A(\adder/adder3/n62 ), .ZN(\adder/g2 ) );
  INV_X1 \adder/adder3/U5  ( .A(\adder/adder3/n101 ), .ZN(\adder/adder3/n60 )
         );
  AOI21_X1 \adder/adder3/U4  ( .B1(\adder/adder3/n64 ), .B2(\adder/adder3/n60 ), .A(SYNOPSYS_UNCONNECTED_42), .ZN(\adder/adder3/n61 ) );
  CLKBUF_X1 \adder/adder3/U3  ( .A(\adder/adder3/n64 ), .Z(\adder/adder3/n56 )
         );
  NOR2_X1 \adder/adder3/U2  ( .A1(alu_operand[17]), .A2(n_2_net__17_), .ZN(
        \adder/adder3/n83 ) );
  OAI21_X2 \adder/adder3/U1  ( .B1(\adder/adder3/n103 ), .B2(
        \adder/adder3/n101 ), .A(\adder/adder3/n77 ), .ZN(\adder/adder3/n106 )
         );
  OAI21_X1 \adder/adder4/U79  ( .B1(\adder/adder4/n61 ), .B2(
        \adder/adder4/n110 ), .A(\adder/adder4/n108 ), .ZN(adder_out[31]) );
  INV_X1 \adder/adder4/U78  ( .A(\adder/adder4/n69 ), .ZN(\adder/adder4/n111 )
         );
  OAI22_X1 \adder/adder4/U77  ( .A1(\adder/adder4/n111 ), .A2(
        \adder/adder4/n92 ), .B1(\adder/adder4/n91 ), .B2(\adder/adder4/n69 ), 
        .ZN(adder_out[26]) );
  XNOR2_X1 \adder/adder4/U76  ( .A(\adder/adder4/n80 ), .B(\adder/adder4/n76 ), 
        .ZN(\adder/overflow ) );
  AOI21_X1 \adder/adder4/U75  ( .B1(\adder/adder4/n76 ), .B2(
        SYNOPSYS_UNCONNECTED_1), .A(SYNOPSYS_UNCONNECTED_33), .ZN(
        \adder/adder4/n80 ) );
  OAI21_X1 \adder/adder4/U74  ( .B1(\adder/adder4/n75 ), .B2(
        \adder/adder4/n104 ), .A(\adder/adder4/n79 ), .ZN(\adder/adder4/n109 )
         );
  OAI21_X1 \adder/adder4/U73  ( .B1(SYNOPSYS_UNCONNECTED_36), .B2(
        \adder/adder4/n96 ), .A(\adder/adder4/n67 ), .ZN(\adder/adder4/n97 )
         );
  OAI21_X1 \adder/adder4/U72  ( .B1(\adder/adder4/n99 ), .B2(
        \adder/adder4/n67 ), .A(\adder/adder4/n97 ), .ZN(adder_out[28]) );
  XNOR2_X1 \adder/adder4/U71  ( .A(\adder/adder4/n106 ), .B(
        \adder/adder4/n105 ), .ZN(adder_out[30]) );
  AOI21_X1 \adder/adder4/U70  ( .B1(\adder/n14 ), .B2(SYNOPSYS_UNCONNECTED_8), 
        .A(SYNOPSYS_UNCONNECTED_40), .ZN(\adder/adder4/n88 ) );
  OAI21_X1 \adder/adder4/U69  ( .B1(\adder/adder4/n88 ), .B2(
        \adder/adder4/n86 ), .A(\adder/adder4/n77 ), .ZN(\adder/adder4/n90 )
         );
  OAI21_X1 \adder/adder4/U68  ( .B1(\adder/adder4/n95 ), .B2(
        \adder/adder4/n93 ), .A(\adder/adder4/n78 ), .ZN(\adder/adder4/n98 )
         );
  XNOR2_X1 \adder/adder4/U67  ( .A(\adder/adder4/n70 ), .B(\adder/adder4/n87 ), 
        .ZN(adder_out[25]) );
  XNOR2_X1 \adder/adder4/U66  ( .A(\adder/adder4/n74 ), .B(\adder/adder4/n94 ), 
        .ZN(adder_out[27]) );
  AOI21_X1 \adder/adder4/U65  ( .B1(\adder/adder4/n90 ), .B2(
        SYNOPSYS_UNCONNECTED_6), .A(SYNOPSYS_UNCONNECTED_38), .ZN(
        \adder/adder4/n95 ) );
  OAI22_X1 \adder/adder4/U64  ( .A1(\adder/adder4/n103 ), .A2(
        \adder/adder4/n72 ), .B1(\adder/adder4/n71 ), .B2(\adder/adder4/n101 ), 
        .ZN(adder_out[29]) );
  CLKBUF_X1 \adder/adder4/U63  ( .A(\adder/adder4/n61 ), .Z(\adder/adder4/n76 ) );
  OAI21_X1 \adder/adder4/U62  ( .B1(SYNOPSYS_UNCONNECTED_40), .B2(
        \adder/adder4/n83 ), .A(\adder/adder4/n64 ), .ZN(\adder/adder4/n84 )
         );
  OAI21_X1 \adder/adder4/U61  ( .B1(\adder/adder4/n85 ), .B2(
        \adder/adder4/n64 ), .A(\adder/adder4/n84 ), .ZN(adder_out[24]) );
  AND2_X1 \adder/adder4/U60  ( .A1(alu_operand[24]), .A2(n_2_net__24_), .ZN(
        SYNOPSYS_UNCONNECTED_40) );
  AND2_X1 \adder/adder4/U59  ( .A1(alu_operand[28]), .A2(n_2_net__28_), .ZN(
        SYNOPSYS_UNCONNECTED_36) );
  AND2_X1 \adder/adder4/U58  ( .A1(n_2_net__31_), .A2(alu_operand[31]), .ZN(
        SYNOPSYS_UNCONNECTED_33) );
  AND2_X1 \adder/adder4/U57  ( .A1(alu_operand[26]), .A2(n_2_net__26_), .ZN(
        SYNOPSYS_UNCONNECTED_38) );
  AND2_X1 \adder/adder4/U56  ( .A1(alu_operand[29]), .A2(n_2_net__29_), .ZN(
        SYNOPSYS_UNCONNECTED_35) );
  NAND2_X1 \adder/adder4/U55  ( .A1(alu_operand[27]), .A2(n_2_net__27_), .ZN(
        \adder/adder4/n78 ) );
  NAND2_X1 \adder/adder4/U54  ( .A1(alu_operand[30]), .A2(n_2_net__30_), .ZN(
        \adder/adder4/n79 ) );
  NAND2_X1 \adder/adder4/U53  ( .A1(alu_operand[25]), .A2(n_2_net__25_), .ZN(
        \adder/adder4/n77 ) );
  NOR2_X1 \adder/adder4/U52  ( .A1(alu_operand[31]), .A2(n_2_net__31_), .ZN(
        \adder/adder4/n107 ) );
  NOR2_X1 \adder/adder4/U51  ( .A1(alu_operand[28]), .A2(n_2_net__28_), .ZN(
        \adder/adder4/n96 ) );
  NOR2_X1 \adder/adder4/U50  ( .A1(alu_operand[24]), .A2(n_2_net__24_), .ZN(
        \adder/adder4/n83 ) );
  NOR2_X1 \adder/adder4/U49  ( .A1(alu_operand[26]), .A2(n_2_net__26_), .ZN(
        \adder/adder4/n89 ) );
  NOR2_X1 \adder/adder4/U48  ( .A1(alu_operand[29]), .A2(n_2_net__29_), .ZN(
        \adder/adder4/n100 ) );
  NOR2_X1 \adder/adder4/U47  ( .A1(alu_operand[27]), .A2(n_2_net__27_), .ZN(
        \adder/adder4/n93 ) );
  NOR2_X1 \adder/adder4/U46  ( .A1(alu_operand[30]), .A2(n_2_net__30_), .ZN(
        \adder/adder4/n104 ) );
  NOR2_X1 \adder/adder4/U45  ( .A1(alu_operand[25]), .A2(n_2_net__25_), .ZN(
        \adder/adder4/n86 ) );
  XNOR2_X1 \adder/adder4/U44  ( .A(n_2_net__31_), .B(alu_operand[31]), .ZN(
        \adder/adder4/n110 ) );
  XNOR2_X1 \adder/adder4/U43  ( .A(n_2_net__24_), .B(alu_operand[24]), .ZN(
        \adder/adder4/n85 ) );
  XNOR2_X1 \adder/adder4/U42  ( .A(n_2_net__28_), .B(alu_operand[28]), .ZN(
        \adder/adder4/n99 ) );
  NOR2_X1 \adder/adder4/U41  ( .A1(SYNOPSYS_UNCONNECTED_35), .A2(
        \adder/adder4/n100 ), .ZN(\adder/adder4/n101 ) );
  XNOR2_X1 \adder/adder4/U40  ( .A(n_2_net__29_), .B(alu_operand[29]), .ZN(
        \adder/adder4/n103 ) );
  NOR2_X1 \adder/adder4/U39  ( .A1(SYNOPSYS_UNCONNECTED_38), .A2(
        \adder/adder4/n89 ), .ZN(\adder/adder4/n92 ) );
  XNOR2_X1 \adder/adder4/U38  ( .A(n_2_net__26_), .B(alu_operand[26]), .ZN(
        \adder/adder4/n91 ) );
  INV_X1 \adder/adder4/U37  ( .A(\adder/adder4/n79 ), .ZN(
        SYNOPSYS_UNCONNECTED_34) );
  INV_X1 \adder/adder4/U36  ( .A(\adder/adder4/n78 ), .ZN(
        SYNOPSYS_UNCONNECTED_37) );
  INV_X1 \adder/adder4/U35  ( .A(\adder/adder4/n77 ), .ZN(
        SYNOPSYS_UNCONNECTED_39) );
  INV_X1 \adder/adder4/U34  ( .A(\adder/adder4/n107 ), .ZN(
        SYNOPSYS_UNCONNECTED_1) );
  INV_X1 \adder/adder4/U33  ( .A(\adder/adder4/n96 ), .ZN(
        SYNOPSYS_UNCONNECTED_4) );
  INV_X1 \adder/adder4/U32  ( .A(\adder/adder4/n83 ), .ZN(
        SYNOPSYS_UNCONNECTED_8) );
  INV_X1 \adder/adder4/U31  ( .A(\adder/adder4/n89 ), .ZN(
        SYNOPSYS_UNCONNECTED_6) );
  INV_X1 \adder/adder4/U30  ( .A(\adder/adder4/n100 ), .ZN(
        SYNOPSYS_UNCONNECTED_3) );
  INV_X1 \adder/adder4/U29  ( .A(\adder/adder4/n86 ), .ZN(
        SYNOPSYS_UNCONNECTED_7) );
  INV_X1 \adder/adder4/U28  ( .A(\adder/adder4/n104 ), .ZN(
        SYNOPSYS_UNCONNECTED_2) );
  INV_X1 \adder/adder4/U27  ( .A(\adder/adder4/n93 ), .ZN(
        SYNOPSYS_UNCONNECTED_5) );
  NAND4_X1 \adder/adder4/U26  ( .A1(SYNOPSYS_UNCONNECTED_5), .A2(
        SYNOPSYS_UNCONNECTED_4), .A3(SYNOPSYS_UNCONNECTED_3), .A4(
        SYNOPSYS_UNCONNECTED_2), .ZN(\adder/adder4/n82 ) );
  NAND4_X1 \adder/adder4/U25  ( .A1(SYNOPSYS_UNCONNECTED_1), .A2(
        SYNOPSYS_UNCONNECTED_8), .A3(SYNOPSYS_UNCONNECTED_7), .A4(
        SYNOPSYS_UNCONNECTED_6), .ZN(\adder/adder4/n81 ) );
  AOI21_X1 \adder/adder4/U24  ( .B1(\adder/adder4/n60 ), .B2(
        SYNOPSYS_UNCONNECTED_3), .A(SYNOPSYS_UNCONNECTED_35), .ZN(
        \adder/adder4/n106 ) );
  NOR2_X1 \adder/adder4/U23  ( .A1(SYNOPSYS_UNCONNECTED_34), .A2(
        \adder/adder4/n104 ), .ZN(\adder/adder4/n105 ) );
  NOR2_X1 \adder/adder4/U22  ( .A1(SYNOPSYS_UNCONNECTED_39), .A2(
        \adder/adder4/n86 ), .ZN(\adder/adder4/n87 ) );
  NOR2_X1 \adder/adder4/U21  ( .A1(SYNOPSYS_UNCONNECTED_37), .A2(
        \adder/adder4/n93 ), .ZN(\adder/adder4/n94 ) );
  INV_X1 \adder/adder4/U20  ( .A(\adder/adder4/n80 ), .ZN(\adder/adder4/gen )
         );
  NOR2_X1 \adder/adder4/U19  ( .A1(\adder/adder4/n82 ), .A2(\adder/adder4/n81 ), .ZN(\adder/adder4/prop ) );
  AOI21_X1 \adder/adder4/U18  ( .B1(\adder/adder4/n69 ), .B2(
        SYNOPSYS_UNCONNECTED_6), .A(SYNOPSYS_UNCONNECTED_38), .ZN(
        \adder/adder4/n74 ) );
  NAND2_X1 \adder/adder4/U17  ( .A1(\adder/adder4/n109 ), .A2(
        \adder/adder4/n73 ), .ZN(\adder/adder4/n108 ) );
  OR2_X1 \adder/adder4/U16  ( .A1(SYNOPSYS_UNCONNECTED_33), .A2(
        \adder/adder4/n107 ), .ZN(\adder/adder4/n73 ) );
  INV_X1 \adder/adder4/U15  ( .A(\adder/adder4/n68 ), .ZN(\adder/adder4/n72 )
         );
  AOI21_X1 \adder/adder4/U14  ( .B1(\adder/adder4/n98 ), .B2(
        SYNOPSYS_UNCONNECTED_4), .A(SYNOPSYS_UNCONNECTED_36), .ZN(
        \adder/adder4/n102 ) );
  INV_X1 \adder/adder4/U13  ( .A(\adder/adder4/n72 ), .ZN(\adder/adder4/n71 )
         );
  AOI21_X1 \adder/adder4/U12  ( .B1(\adder/adder4/n64 ), .B2(
        SYNOPSYS_UNCONNECTED_8), .A(SYNOPSYS_UNCONNECTED_40), .ZN(
        \adder/adder4/n70 ) );
  CLKBUF_X1 \adder/adder4/U11  ( .A(\adder/adder4/n65 ), .Z(\adder/adder4/n69 ) );
  AOI21_X1 \adder/adder4/U10  ( .B1(\adder/adder4/n67 ), .B2(
        SYNOPSYS_UNCONNECTED_4), .A(SYNOPSYS_UNCONNECTED_36), .ZN(
        \adder/adder4/n68 ) );
  OAI21_X1 \adder/adder4/U9  ( .B1(\adder/adder4/n66 ), .B2(\adder/adder4/n93 ), .A(\adder/adder4/n78 ), .ZN(\adder/adder4/n67 ) );
  AOI21_X1 \adder/adder4/U8  ( .B1(\adder/adder4/n65 ), .B2(
        SYNOPSYS_UNCONNECTED_6), .A(SYNOPSYS_UNCONNECTED_38), .ZN(
        \adder/adder4/n66 ) );
  CLKBUF_X1 \adder/adder4/U7  ( .A(\adder/adder4/n90 ), .Z(\adder/adder4/n65 )
         );
  CLKBUF_X1 \adder/adder4/U6  ( .A(\adder/n14 ), .Z(\adder/adder4/n64 ) );
  INV_X1 \adder/adder4/U5  ( .A(\adder/adder4/n63 ), .ZN(\adder/adder4/n75 )
         );
  INV_X1 \adder/adder4/U4  ( .A(SYNOPSYS_UNCONNECTED_35), .ZN(
        \adder/adder4/n62 ) );
  OAI21_X1 \adder/adder4/U3  ( .B1(\adder/adder4/n102 ), .B2(
        \adder/adder4/n100 ), .A(\adder/adder4/n62 ), .ZN(\adder/adder4/n63 )
         );
  OAI21_X1 \adder/adder4/U2  ( .B1(\adder/adder4/n75 ), .B2(
        \adder/adder4/n104 ), .A(\adder/adder4/n79 ), .ZN(\adder/adder4/n61 )
         );
  CLKBUF_X1 \adder/adder4/U1  ( .A(\adder/adder4/n72 ), .Z(\adder/adder4/n60 )
         );
  AOI21_X1 \adder_sign/U8  ( .B1(\adder_sign/p2 ), .B2(\adder_sign/n16 ), .A(
        \adder_sign/g2 ), .ZN(\adder_sign/n14 ) );
  INV_X1 \adder_sign/U7  ( .A(\adder_sign/n14 ), .ZN(\adder_sign/n17 ) );
  AND2_X1 \adder_sign/U6  ( .A1(\adder_sign/n15 ), .A2(\adder_sign/p1 ), .ZN(
        \adder_sign/n13 ) );
  OR2_X2 \adder_sign/U5  ( .A1(\adder_sign/n13 ), .A2(\adder_sign/g1 ), .ZN(
        \adder_sign/n16 ) );
  INV_X1 \adder_sign/U4  ( .A(\adder_sign/g0 ), .ZN(\adder_sign/n12 ) );
  INV_X1 \adder_sign/U3  ( .A(1'b0), .ZN(\adder_sign/n11 ) );
  INV_X1 \adder_sign/U2  ( .A(\adder_sign/p0 ), .ZN(\adder_sign/n10 ) );
  OAI21_X1 \adder_sign/U1  ( .B1(\adder_sign/n10 ), .B2(\adder_sign/n11 ), .A(
        \adder_sign/n12 ), .ZN(\adder_sign/n15 ) );
  NOR2_X1 \adder_sign/adder1/U71  ( .A1(1'b1), .A2(n579), .ZN(
        \adder_sign/adder1/n74 ) );
  AND2_X1 \adder_sign/adder1/U70  ( .A1(1'b1), .A2(n579), .ZN(
        SYNOPSYS_UNCONNECTED_128) );
  XNOR2_X1 \adder_sign/adder1/U69  ( .A(n579), .B(1'b1), .ZN(
        \adder_sign/adder1/n76 ) );
  AND2_X1 \adder_sign/adder1/U68  ( .A1(1'b0), .A2(n583), .ZN(
        SYNOPSYS_UNCONNECTED_124) );
  AND2_X1 \adder_sign/adder1/U67  ( .A1(1'b0), .A2(n584), .ZN(
        SYNOPSYS_UNCONNECTED_123) );
  AND2_X1 \adder_sign/adder1/U66  ( .A1(1'b0), .A2(n581), .ZN(
        SYNOPSYS_UNCONNECTED_126) );
  AND2_X1 \adder_sign/adder1/U65  ( .A1(n586), .A2(1'b0), .ZN(
        SYNOPSYS_UNCONNECTED_121) );
  NAND2_X1 \adder_sign/adder1/U64  ( .A1(1'b0), .A2(n585), .ZN(
        \adder_sign/adder1/n70 ) );
  NAND2_X1 \adder_sign/adder1/U63  ( .A1(1'b0), .A2(n582), .ZN(
        \adder_sign/adder1/n69 ) );
  NAND2_X1 \adder_sign/adder1/U62  ( .A1(1'b0), .A2(n580), .ZN(
        \adder_sign/adder1/n68 ) );
  NOR2_X1 \adder_sign/adder1/U61  ( .A1(SYNOPSYS_UNCONNECTED_123), .A2(
        \adder_sign/adder1/n91 ), .ZN(\adder_sign/adder1/n92 ) );
  XNOR2_X1 \adder_sign/adder1/U60  ( .A(n584), .B(1'b0), .ZN(
        \adder_sign/adder1/n94 ) );
  OAI22_X1 \adder_sign/adder1/U59  ( .A1(\adder_sign/adder1/n94 ), .A2(
        \adder_sign/adder1/n104 ), .B1(\adder_sign/adder1/n66 ), .B2(
        \adder_sign/adder1/n92 ), .ZN(sign_fixed[5]) );
  OAI21_X1 \adder_sign/adder1/U58  ( .B1(SYNOPSYS_UNCONNECTED_121), .B2(
        \adder_sign/adder1/n98 ), .A(\adder_sign/adder1/n60 ), .ZN(
        \adder_sign/adder1/n99 ) );
  XNOR2_X1 \adder_sign/adder1/U57  ( .A(n586), .B(1'b0), .ZN(
        \adder_sign/adder1/n101 ) );
  OAI21_X1 \adder_sign/adder1/U56  ( .B1(\adder_sign/adder1/n101 ), .B2(
        \adder_sign/adder1/n60 ), .A(\adder_sign/adder1/n99 ), .ZN(
        sign_fixed[7]) );
  OAI21_X1 \adder_sign/adder1/U55  ( .B1(SYNOPSYS_UNCONNECTED_128), .B2(
        \adder_sign/adder1/n74 ), .A(1'b0), .ZN(\adder_sign/adder1/n75 ) );
  OAI21_X1 \adder_sign/adder1/U54  ( .B1(1'b0), .B2(\adder_sign/adder1/n76 ), 
        .A(\adder_sign/adder1/n75 ), .ZN(sign_fixed[0]) );
  OAI21_X1 \adder_sign/adder1/U53  ( .B1(SYNOPSYS_UNCONNECTED_124), .B2(
        \adder_sign/adder1/n87 ), .A(\adder_sign/adder1/n67 ), .ZN(
        \adder_sign/adder1/n88 ) );
  XNOR2_X1 \adder_sign/adder1/U52  ( .A(n583), .B(1'b0), .ZN(
        \adder_sign/adder1/n90 ) );
  OAI21_X1 \adder_sign/adder1/U51  ( .B1(\adder_sign/adder1/n90 ), .B2(
        \adder_sign/adder1/n67 ), .A(\adder_sign/adder1/n88 ), .ZN(
        sign_fixed[4]) );
  INV_X1 \adder_sign/adder1/U50  ( .A(\adder_sign/adder1/n64 ), .ZN(
        \adder_sign/adder1/n103 ) );
  NOR2_X1 \adder_sign/adder1/U49  ( .A1(SYNOPSYS_UNCONNECTED_126), .A2(
        \adder_sign/adder1/n80 ), .ZN(\adder_sign/adder1/n83 ) );
  XNOR2_X1 \adder_sign/adder1/U48  ( .A(n581), .B(1'b0), .ZN(
        \adder_sign/adder1/n82 ) );
  OAI22_X1 \adder_sign/adder1/U47  ( .A1(\adder_sign/adder1/n103 ), .A2(
        \adder_sign/adder1/n83 ), .B1(\adder_sign/adder1/n82 ), .B2(
        \adder_sign/adder1/n64 ), .ZN(sign_fixed[2]) );
  NOR2_X1 \adder_sign/adder1/U46  ( .A1(\adder_sign/adder1/n73 ), .A2(
        \adder_sign/adder1/n72 ), .ZN(\adder_sign/p0 ) );
  AOI21_X1 \adder_sign/adder1/U45  ( .B1(SYNOPSYS_UNCONNECTED_96), .B2(1'b0), 
        .A(SYNOPSYS_UNCONNECTED_128), .ZN(\adder_sign/adder1/n79 ) );
  NOR2_X1 \adder_sign/adder1/U44  ( .A1(1'b0), .A2(n586), .ZN(
        \adder_sign/adder1/n98 ) );
  NOR2_X1 \adder_sign/adder1/U43  ( .A1(1'b0), .A2(n583), .ZN(
        \adder_sign/adder1/n87 ) );
  NOR2_X1 \adder_sign/adder1/U42  ( .A1(1'b0), .A2(n581), .ZN(
        \adder_sign/adder1/n80 ) );
  NOR2_X1 \adder_sign/adder1/U41  ( .A1(1'b0), .A2(n584), .ZN(
        \adder_sign/adder1/n91 ) );
  NOR2_X1 \adder_sign/adder1/U40  ( .A1(1'b0), .A2(n582), .ZN(
        \adder_sign/adder1/n84 ) );
  NOR2_X1 \adder_sign/adder1/U39  ( .A1(1'b0), .A2(n585), .ZN(
        \adder_sign/adder1/n95 ) );
  INV_X1 \adder_sign/adder1/U38  ( .A(\adder_sign/adder1/n70 ), .ZN(
        SYNOPSYS_UNCONNECTED_122) );
  INV_X1 \adder_sign/adder1/U37  ( .A(\adder_sign/adder1/n69 ), .ZN(
        SYNOPSYS_UNCONNECTED_125) );
  INV_X1 \adder_sign/adder1/U36  ( .A(\adder_sign/adder1/n68 ), .ZN(
        SYNOPSYS_UNCONNECTED_127) );
  INV_X1 \adder_sign/adder1/U35  ( .A(\adder_sign/adder1/n98 ), .ZN(
        SYNOPSYS_UNCONNECTED_89) );
  INV_X1 \adder_sign/adder1/U34  ( .A(\adder_sign/adder1/n87 ), .ZN(
        SYNOPSYS_UNCONNECTED_92) );
  INV_X1 \adder_sign/adder1/U33  ( .A(\adder_sign/adder1/n91 ), .ZN(
        SYNOPSYS_UNCONNECTED_91) );
  INV_X1 \adder_sign/adder1/U32  ( .A(\adder_sign/adder1/n80 ), .ZN(
        SYNOPSYS_UNCONNECTED_94) );
  INV_X1 \adder_sign/adder1/U31  ( .A(\adder_sign/adder1/n95 ), .ZN(
        SYNOPSYS_UNCONNECTED_90) );
  INV_X1 \adder_sign/adder1/U30  ( .A(\adder_sign/adder1/n84 ), .ZN(
        SYNOPSYS_UNCONNECTED_93) );
  INV_X1 \adder_sign/adder1/U29  ( .A(\adder_sign/adder1/n77 ), .ZN(
        SYNOPSYS_UNCONNECTED_95) );
  INV_X1 \adder_sign/adder1/U28  ( .A(\adder_sign/adder1/n74 ), .ZN(
        SYNOPSYS_UNCONNECTED_96) );
  NAND4_X1 \adder_sign/adder1/U27  ( .A1(SYNOPSYS_UNCONNECTED_93), .A2(
        SYNOPSYS_UNCONNECTED_92), .A3(SYNOPSYS_UNCONNECTED_91), .A4(
        SYNOPSYS_UNCONNECTED_90), .ZN(\adder_sign/adder1/n73 ) );
  NAND4_X1 \adder_sign/adder1/U26  ( .A1(SYNOPSYS_UNCONNECTED_89), .A2(
        SYNOPSYS_UNCONNECTED_96), .A3(SYNOPSYS_UNCONNECTED_95), .A4(
        SYNOPSYS_UNCONNECTED_94), .ZN(\adder_sign/adder1/n72 ) );
  NOR2_X1 \adder_sign/adder1/U25  ( .A1(SYNOPSYS_UNCONNECTED_122), .A2(
        \adder_sign/adder1/n95 ), .ZN(\adder_sign/adder1/n96 ) );
  XNOR2_X1 \adder_sign/adder1/U24  ( .A(\adder_sign/adder1/n65 ), .B(
        \adder_sign/adder1/n96 ), .ZN(sign_fixed[6]) );
  NOR2_X1 \adder_sign/adder1/U23  ( .A1(SYNOPSYS_UNCONNECTED_127), .A2(
        \adder_sign/adder1/n77 ), .ZN(\adder_sign/adder1/n78 ) );
  XNOR2_X1 \adder_sign/adder1/U22  ( .A(\adder_sign/adder1/n79 ), .B(
        \adder_sign/adder1/n78 ), .ZN(sign_fixed[1]) );
  NOR2_X1 \adder_sign/adder1/U21  ( .A1(SYNOPSYS_UNCONNECTED_125), .A2(
        \adder_sign/adder1/n84 ), .ZN(\adder_sign/adder1/n85 ) );
  XNOR2_X1 \adder_sign/adder1/U20  ( .A(\adder_sign/adder1/n86 ), .B(
        \adder_sign/adder1/n85 ), .ZN(sign_fixed[3]) );
  AOI21_X1 \adder_sign/adder1/U19  ( .B1(\adder_sign/adder1/n89 ), .B2(
        SYNOPSYS_UNCONNECTED_92), .A(SYNOPSYS_UNCONNECTED_124), .ZN(
        \adder_sign/adder1/n93 ) );
  AOI21_X1 \adder_sign/adder1/U18  ( .B1(\adder_sign/adder1/n81 ), .B2(
        SYNOPSYS_UNCONNECTED_94), .A(SYNOPSYS_UNCONNECTED_126), .ZN(
        \adder_sign/adder1/n86 ) );
  AOI21_X1 \adder_sign/adder1/U17  ( .B1(\adder_sign/adder1/n60 ), .B2(
        SYNOPSYS_UNCONNECTED_89), .A(SYNOPSYS_UNCONNECTED_121), .ZN(
        \adder_sign/adder1/n71 ) );
  OAI21_X1 \adder_sign/adder1/U16  ( .B1(\adder_sign/adder1/n86 ), .B2(
        \adder_sign/adder1/n84 ), .A(\adder_sign/adder1/n69 ), .ZN(
        \adder_sign/adder1/n89 ) );
  OAI21_X1 \adder_sign/adder1/U15  ( .B1(\adder_sign/adder1/n79 ), .B2(
        \adder_sign/adder1/n77 ), .A(\adder_sign/adder1/n68 ), .ZN(
        \adder_sign/adder1/n81 ) );
  XNOR2_X1 \adder_sign/adder1/U14  ( .A(\adder_sign/adder1/n71 ), .B(
        \adder_sign/adder1/n60 ), .ZN(\adder_sign/adder1/overflow ) );
  INV_X1 \adder_sign/adder1/U13  ( .A(\adder_sign/adder1/n93 ), .ZN(
        \adder_sign/adder1/n104 ) );
  CLKBUF_X1 \adder_sign/adder1/U12  ( .A(\adder_sign/adder1/n89 ), .Z(
        \adder_sign/adder1/n67 ) );
  INV_X1 \adder_sign/adder1/U11  ( .A(\adder_sign/adder1/n104 ), .ZN(
        \adder_sign/adder1/n66 ) );
  AOI21_X1 \adder_sign/adder1/U10  ( .B1(\adder_sign/adder1/n104 ), .B2(
        SYNOPSYS_UNCONNECTED_91), .A(SYNOPSYS_UNCONNECTED_123), .ZN(
        \adder_sign/adder1/n65 ) );
  NOR2_X1 \adder_sign/adder1/U9  ( .A1(1'b0), .A2(n580), .ZN(
        \adder_sign/adder1/n77 ) );
  CLKBUF_X1 \adder_sign/adder1/U8  ( .A(\adder_sign/adder1/n81 ), .Z(
        \adder_sign/adder1/n64 ) );
  INV_X1 \adder_sign/adder1/U7  ( .A(\adder_sign/adder1/n63 ), .ZN(
        \adder_sign/adder1/n97 ) );
  INV_X1 \adder_sign/adder1/U6  ( .A(SYNOPSYS_UNCONNECTED_123), .ZN(
        \adder_sign/adder1/n62 ) );
  OAI21_X1 \adder_sign/adder1/U5  ( .B1(\adder_sign/adder1/n91 ), .B2(
        \adder_sign/adder1/n93 ), .A(\adder_sign/adder1/n62 ), .ZN(
        \adder_sign/adder1/n63 ) );
  INV_X1 \adder_sign/adder1/U4  ( .A(\adder_sign/adder1/n61 ), .ZN(
        \adder_sign/g0 ) );
  AOI21_X1 \adder_sign/adder1/U3  ( .B1(SYNOPSYS_UNCONNECTED_89), .B2(
        \adder_sign/adder1/n100 ), .A(SYNOPSYS_UNCONNECTED_121), .ZN(
        \adder_sign/adder1/n61 ) );
  OAI21_X1 \adder_sign/adder1/U2  ( .B1(\adder_sign/adder1/n97 ), .B2(
        \adder_sign/adder1/n95 ), .A(\adder_sign/adder1/n70 ), .ZN(
        \adder_sign/adder1/n100 ) );
  CLKBUF_X1 \adder_sign/adder1/U1  ( .A(\adder_sign/adder1/n100 ), .Z(
        \adder_sign/adder1/n60 ) );
  AND2_X1 \adder_sign/adder2/U73  ( .A1(1'b0), .A2(n587), .ZN(
        SYNOPSYS_UNCONNECTED_120) );
  AND2_X1 \adder_sign/adder2/U72  ( .A1(1'b0), .A2(n591), .ZN(
        SYNOPSYS_UNCONNECTED_116) );
  AND2_X1 \adder_sign/adder2/U71  ( .A1(1'b0), .A2(n589), .ZN(
        SYNOPSYS_UNCONNECTED_118) );
  AND2_X1 \adder_sign/adder2/U70  ( .A1(1'b0), .A2(n592), .ZN(
        SYNOPSYS_UNCONNECTED_115) );
  AND2_X1 \adder_sign/adder2/U69  ( .A1(n594), .A2(1'b0), .ZN(
        SYNOPSYS_UNCONNECTED_113) );
  NAND2_X1 \adder_sign/adder2/U68  ( .A1(1'b0), .A2(n593), .ZN(
        \adder_sign/adder2/n72 ) );
  NAND2_X1 \adder_sign/adder2/U67  ( .A1(1'b0), .A2(n590), .ZN(
        \adder_sign/adder2/n71 ) );
  NAND2_X1 \adder_sign/adder2/U66  ( .A1(1'b0), .A2(n588), .ZN(
        \adder_sign/adder2/n70 ) );
  OAI21_X1 \adder_sign/adder2/U65  ( .B1(SYNOPSYS_UNCONNECTED_120), .B2(
        \adder_sign/adder2/n76 ), .A(\adder_sign/n15 ), .ZN(
        \adder_sign/adder2/n77 ) );
  XNOR2_X1 \adder_sign/adder2/U64  ( .A(n587), .B(1'b0), .ZN(
        \adder_sign/adder2/n78 ) );
  OAI21_X1 \adder_sign/adder2/U63  ( .B1(\adder_sign/n15 ), .B2(
        \adder_sign/adder2/n78 ), .A(\adder_sign/adder2/n77 ), .ZN(
        sign_fixed[8]) );
  OAI21_X1 \adder_sign/adder2/U62  ( .B1(SYNOPSYS_UNCONNECTED_116), .B2(
        \adder_sign/adder2/n89 ), .A(\adder_sign/adder2/n60 ), .ZN(
        \adder_sign/adder2/n90 ) );
  XNOR2_X1 \adder_sign/adder2/U61  ( .A(n591), .B(1'b0), .ZN(
        \adder_sign/adder2/n92 ) );
  OAI21_X1 \adder_sign/adder2/U60  ( .B1(\adder_sign/adder2/n92 ), .B2(
        \adder_sign/adder2/n60 ), .A(\adder_sign/adder2/n90 ), .ZN(
        sign_fixed[12]) );
  OAI21_X1 \adder_sign/adder2/U59  ( .B1(SYNOPSYS_UNCONNECTED_113), .B2(
        \adder_sign/adder2/n100 ), .A(\adder_sign/adder2/n62 ), .ZN(
        \adder_sign/adder2/n101 ) );
  XNOR2_X1 \adder_sign/adder2/U58  ( .A(n594), .B(1'b0), .ZN(
        \adder_sign/adder2/n103 ) );
  OAI21_X1 \adder_sign/adder2/U57  ( .B1(\adder_sign/adder2/n103 ), .B2(
        \adder_sign/adder2/n62 ), .A(\adder_sign/adder2/n101 ), .ZN(
        sign_fixed[15]) );
  NOR2_X1 \adder_sign/adder2/U56  ( .A1(1'b0), .A2(n594), .ZN(
        \adder_sign/adder2/n100 ) );
  NOR2_X1 \adder_sign/adder2/U55  ( .A1(1'b0), .A2(n591), .ZN(
        \adder_sign/adder2/n89 ) );
  NOR2_X1 \adder_sign/adder2/U54  ( .A1(1'b0), .A2(n589), .ZN(
        \adder_sign/adder2/n82 ) );
  NOR2_X1 \adder_sign/adder2/U53  ( .A1(SYNOPSYS_UNCONNECTED_115), .A2(
        \adder_sign/adder2/n93 ), .ZN(\adder_sign/adder2/n94 ) );
  XNOR2_X1 \adder_sign/adder2/U52  ( .A(n592), .B(1'b0), .ZN(
        \adder_sign/adder2/n96 ) );
  OAI22_X1 \adder_sign/adder2/U51  ( .A1(\adder_sign/adder2/n96 ), .A2(
        \adder_sign/adder2/n105 ), .B1(\adder_sign/adder2/n69 ), .B2(
        \adder_sign/adder2/n94 ), .ZN(sign_fixed[13]) );
  INV_X1 \adder_sign/adder2/U50  ( .A(\adder_sign/adder2/n61 ), .ZN(
        \adder_sign/adder2/n104 ) );
  NOR2_X1 \adder_sign/adder2/U49  ( .A1(SYNOPSYS_UNCONNECTED_118), .A2(
        \adder_sign/adder2/n82 ), .ZN(\adder_sign/adder2/n85 ) );
  XNOR2_X1 \adder_sign/adder2/U48  ( .A(n589), .B(1'b0), .ZN(
        \adder_sign/adder2/n84 ) );
  OAI22_X1 \adder_sign/adder2/U47  ( .A1(\adder_sign/adder2/n104 ), .A2(
        \adder_sign/adder2/n85 ), .B1(\adder_sign/adder2/n84 ), .B2(
        \adder_sign/adder2/n61 ), .ZN(sign_fixed[10]) );
  NOR2_X1 \adder_sign/adder2/U46  ( .A1(1'b0), .A2(n593), .ZN(
        \adder_sign/adder2/n97 ) );
  NOR2_X1 \adder_sign/adder2/U45  ( .A1(1'b0), .A2(n590), .ZN(
        \adder_sign/adder2/n86 ) );
  NOR2_X1 \adder_sign/adder2/U44  ( .A1(1'b0), .A2(n588), .ZN(
        \adder_sign/adder2/n79 ) );
  NOR2_X1 \adder_sign/adder2/U43  ( .A1(1'b0), .A2(n587), .ZN(
        \adder_sign/adder2/n76 ) );
  INV_X1 \adder_sign/adder2/U42  ( .A(\adder_sign/adder2/n70 ), .ZN(
        SYNOPSYS_UNCONNECTED_119) );
  INV_X1 \adder_sign/adder2/U41  ( .A(\adder_sign/adder2/n72 ), .ZN(
        SYNOPSYS_UNCONNECTED_114) );
  INV_X1 \adder_sign/adder2/U40  ( .A(\adder_sign/adder2/n71 ), .ZN(
        SYNOPSYS_UNCONNECTED_117) );
  INV_X1 \adder_sign/adder2/U39  ( .A(\adder_sign/adder2/n100 ), .ZN(
        SYNOPSYS_UNCONNECTED_81) );
  INV_X1 \adder_sign/adder2/U38  ( .A(\adder_sign/adder2/n89 ), .ZN(
        SYNOPSYS_UNCONNECTED_84) );
  INV_X1 \adder_sign/adder2/U37  ( .A(\adder_sign/adder2/n93 ), .ZN(
        SYNOPSYS_UNCONNECTED_83) );
  INV_X1 \adder_sign/adder2/U36  ( .A(\adder_sign/adder2/n76 ), .ZN(
        SYNOPSYS_UNCONNECTED_88) );
  INV_X1 \adder_sign/adder2/U35  ( .A(\adder_sign/adder2/n82 ), .ZN(
        SYNOPSYS_UNCONNECTED_86) );
  INV_X1 \adder_sign/adder2/U34  ( .A(\adder_sign/adder2/n97 ), .ZN(
        SYNOPSYS_UNCONNECTED_82) );
  INV_X1 \adder_sign/adder2/U33  ( .A(\adder_sign/adder2/n79 ), .ZN(
        SYNOPSYS_UNCONNECTED_87) );
  INV_X1 \adder_sign/adder2/U32  ( .A(\adder_sign/adder2/n86 ), .ZN(
        SYNOPSYS_UNCONNECTED_85) );
  NOR2_X1 \adder_sign/adder2/U31  ( .A1(SYNOPSYS_UNCONNECTED_119), .A2(
        \adder_sign/adder2/n79 ), .ZN(\adder_sign/adder2/n80 ) );
  XNOR2_X1 \adder_sign/adder2/U30  ( .A(\adder_sign/adder2/n65 ), .B(
        \adder_sign/adder2/n80 ), .ZN(sign_fixed[9]) );
  NAND4_X1 \adder_sign/adder2/U29  ( .A1(SYNOPSYS_UNCONNECTED_85), .A2(
        SYNOPSYS_UNCONNECTED_84), .A3(SYNOPSYS_UNCONNECTED_83), .A4(
        SYNOPSYS_UNCONNECTED_82), .ZN(\adder_sign/adder2/n75 ) );
  NAND4_X1 \adder_sign/adder2/U28  ( .A1(SYNOPSYS_UNCONNECTED_81), .A2(
        SYNOPSYS_UNCONNECTED_88), .A3(SYNOPSYS_UNCONNECTED_87), .A4(
        SYNOPSYS_UNCONNECTED_86), .ZN(\adder_sign/adder2/n74 ) );
  NOR2_X1 \adder_sign/adder2/U27  ( .A1(SYNOPSYS_UNCONNECTED_114), .A2(
        \adder_sign/adder2/n97 ), .ZN(\adder_sign/adder2/n98 ) );
  XNOR2_X1 \adder_sign/adder2/U26  ( .A(\adder_sign/adder2/n68 ), .B(
        \adder_sign/adder2/n98 ), .ZN(sign_fixed[14]) );
  NOR2_X1 \adder_sign/adder2/U25  ( .A1(SYNOPSYS_UNCONNECTED_117), .A2(
        \adder_sign/adder2/n86 ), .ZN(\adder_sign/adder2/n87 ) );
  XNOR2_X1 \adder_sign/adder2/U24  ( .A(\adder_sign/adder2/n67 ), .B(
        \adder_sign/adder2/n87 ), .ZN(sign_fixed[11]) );
  INV_X1 \adder_sign/adder2/U23  ( .A(\adder_sign/adder2/n73 ), .ZN(
        \adder_sign/g1 ) );
  NOR2_X1 \adder_sign/adder2/U22  ( .A1(\adder_sign/adder2/n75 ), .A2(
        \adder_sign/adder2/n74 ), .ZN(\adder_sign/p1 ) );
  AOI21_X1 \adder_sign/adder2/U21  ( .B1(\adder_sign/adder2/n91 ), .B2(
        SYNOPSYS_UNCONNECTED_84), .A(SYNOPSYS_UNCONNECTED_116), .ZN(
        \adder_sign/adder2/n95 ) );
  AOI21_X1 \adder_sign/adder2/U20  ( .B1(SYNOPSYS_UNCONNECTED_88), .B2(
        \adder_sign/n15 ), .A(SYNOPSYS_UNCONNECTED_120), .ZN(
        \adder_sign/adder2/n81 ) );
  AOI21_X1 \adder_sign/adder2/U19  ( .B1(\adder_sign/adder2/n102 ), .B2(
        SYNOPSYS_UNCONNECTED_81), .A(SYNOPSYS_UNCONNECTED_113), .ZN(
        \adder_sign/adder2/n73 ) );
  OAI21_X1 \adder_sign/adder2/U18  ( .B1(\adder_sign/adder2/n88 ), .B2(
        \adder_sign/adder2/n86 ), .A(\adder_sign/adder2/n71 ), .ZN(
        \adder_sign/adder2/n91 ) );
  OAI21_X1 \adder_sign/adder2/U17  ( .B1(\adder_sign/adder2/n81 ), .B2(
        \adder_sign/adder2/n79 ), .A(\adder_sign/adder2/n70 ), .ZN(
        \adder_sign/adder2/n83 ) );
  XNOR2_X1 \adder_sign/adder2/U16  ( .A(\adder_sign/adder2/n66 ), .B(
        \adder_sign/adder2/n62 ), .ZN(\adder_sign/adder2/overflow ) );
  INV_X1 \adder_sign/adder2/U15  ( .A(\adder_sign/adder2/n95 ), .ZN(
        \adder_sign/adder2/n105 ) );
  INV_X1 \adder_sign/adder2/U14  ( .A(\adder_sign/adder2/n105 ), .ZN(
        \adder_sign/adder2/n69 ) );
  CLKBUF_X1 \adder_sign/adder2/U13  ( .A(\adder_sign/adder2/n99 ), .Z(
        \adder_sign/adder2/n68 ) );
  AOI21_X1 \adder_sign/adder2/U12  ( .B1(\adder_sign/adder2/n83 ), .B2(
        SYNOPSYS_UNCONNECTED_86), .A(SYNOPSYS_UNCONNECTED_118), .ZN(
        \adder_sign/adder2/n88 ) );
  AOI21_X1 \adder_sign/adder2/U11  ( .B1(\adder_sign/adder2/n61 ), .B2(
        SYNOPSYS_UNCONNECTED_86), .A(SYNOPSYS_UNCONNECTED_118), .ZN(
        \adder_sign/adder2/n67 ) );
  OAI21_X1 \adder_sign/adder2/U10  ( .B1(\adder_sign/adder2/n99 ), .B2(
        \adder_sign/adder2/n97 ), .A(\adder_sign/adder2/n72 ), .ZN(
        \adder_sign/adder2/n102 ) );
  INV_X1 \adder_sign/adder2/U9  ( .A(\adder_sign/g1 ), .ZN(
        \adder_sign/adder2/n66 ) );
  CLKBUF_X1 \adder_sign/adder2/U8  ( .A(\adder_sign/adder2/n81 ), .Z(
        \adder_sign/adder2/n65 ) );
  INV_X1 \adder_sign/adder2/U7  ( .A(\adder_sign/adder2/n64 ), .ZN(
        \adder_sign/adder2/n99 ) );
  INV_X1 \adder_sign/adder2/U6  ( .A(SYNOPSYS_UNCONNECTED_115), .ZN(
        \adder_sign/adder2/n63 ) );
  OAI21_X1 \adder_sign/adder2/U5  ( .B1(\adder_sign/adder2/n93 ), .B2(
        \adder_sign/adder2/n95 ), .A(\adder_sign/adder2/n63 ), .ZN(
        \adder_sign/adder2/n64 ) );
  CLKBUF_X1 \adder_sign/adder2/U4  ( .A(\adder_sign/adder2/n102 ), .Z(
        \adder_sign/adder2/n62 ) );
  CLKBUF_X1 \adder_sign/adder2/U3  ( .A(\adder_sign/adder2/n83 ), .Z(
        \adder_sign/adder2/n61 ) );
  CLKBUF_X1 \adder_sign/adder2/U2  ( .A(\adder_sign/adder2/n91 ), .Z(
        \adder_sign/adder2/n60 ) );
  NOR2_X1 \adder_sign/adder2/U1  ( .A1(1'b0), .A2(n592), .ZN(
        \adder_sign/adder2/n93 ) );
  AND2_X1 \adder_sign/adder3/U72  ( .A1(1'b0), .A2(n599), .ZN(
        SYNOPSYS_UNCONNECTED_108) );
  AND2_X1 \adder_sign/adder3/U71  ( .A1(1'b0), .A2(n595), .ZN(
        SYNOPSYS_UNCONNECTED_112) );
  AND2_X1 \adder_sign/adder3/U70  ( .A1(1'b0), .A2(n600), .ZN(
        SYNOPSYS_UNCONNECTED_107) );
  AND2_X1 \adder_sign/adder3/U69  ( .A1(1'b0), .A2(n597), .ZN(
        SYNOPSYS_UNCONNECTED_110) );
  AND2_X1 \adder_sign/adder3/U68  ( .A1(n602), .A2(1'b0), .ZN(
        SYNOPSYS_UNCONNECTED_105) );
  NAND2_X1 \adder_sign/adder3/U67  ( .A1(1'b0), .A2(n601), .ZN(
        \adder_sign/adder3/n71 ) );
  NAND2_X1 \adder_sign/adder3/U66  ( .A1(1'b0), .A2(n598), .ZN(
        \adder_sign/adder3/n70 ) );
  NAND2_X1 \adder_sign/adder3/U65  ( .A1(1'b0), .A2(n596), .ZN(
        \adder_sign/adder3/n69 ) );
  NOR2_X1 \adder_sign/adder3/U64  ( .A1(SYNOPSYS_UNCONNECTED_107), .A2(
        \adder_sign/adder3/n92 ), .ZN(\adder_sign/adder3/n93 ) );
  XNOR2_X1 \adder_sign/adder3/U63  ( .A(n600), .B(1'b0), .ZN(
        \adder_sign/adder3/n95 ) );
  OAI22_X1 \adder_sign/adder3/U62  ( .A1(\adder_sign/adder3/n95 ), .A2(
        \adder_sign/adder3/n104 ), .B1(\adder_sign/adder3/n62 ), .B2(
        \adder_sign/adder3/n93 ), .ZN(sign_fixed[21]) );
  OAI21_X1 \adder_sign/adder3/U61  ( .B1(SYNOPSYS_UNCONNECTED_108), .B2(
        \adder_sign/adder3/n88 ), .A(\adder_sign/adder3/n90 ), .ZN(
        \adder_sign/adder3/n89 ) );
  XNOR2_X1 \adder_sign/adder3/U60  ( .A(n599), .B(1'b0), .ZN(
        \adder_sign/adder3/n91 ) );
  OAI21_X1 \adder_sign/adder3/U59  ( .B1(\adder_sign/adder3/n91 ), .B2(
        \adder_sign/adder3/n90 ), .A(\adder_sign/adder3/n89 ), .ZN(
        sign_fixed[20]) );
  OAI21_X1 \adder_sign/adder3/U58  ( .B1(SYNOPSYS_UNCONNECTED_112), .B2(
        \adder_sign/adder3/n75 ), .A(\adder_sign/n16 ), .ZN(
        \adder_sign/adder3/n76 ) );
  XNOR2_X1 \adder_sign/adder3/U57  ( .A(n595), .B(1'b0), .ZN(
        \adder_sign/adder3/n77 ) );
  OAI21_X1 \adder_sign/adder3/U56  ( .B1(\adder_sign/n16 ), .B2(
        \adder_sign/adder3/n77 ), .A(\adder_sign/adder3/n76 ), .ZN(
        sign_fixed[16]) );
  NOR2_X1 \adder_sign/adder3/U55  ( .A1(1'b0), .A2(n602), .ZN(
        \adder_sign/adder3/n99 ) );
  NOR2_X1 \adder_sign/adder3/U54  ( .A1(1'b0), .A2(n599), .ZN(
        \adder_sign/adder3/n88 ) );
  NOR2_X1 \adder_sign/adder3/U53  ( .A1(1'b0), .A2(n595), .ZN(
        \adder_sign/adder3/n75 ) );
  NOR2_X1 \adder_sign/adder3/U52  ( .A1(1'b0), .A2(n597), .ZN(
        \adder_sign/adder3/n81 ) );
  NOR2_X1 \adder_sign/adder3/U51  ( .A1(1'b0), .A2(n600), .ZN(
        \adder_sign/adder3/n92 ) );
  INV_X1 \adder_sign/adder3/U50  ( .A(\adder_sign/adder3/n63 ), .ZN(
        \adder_sign/adder3/n103 ) );
  NOR2_X1 \adder_sign/adder3/U49  ( .A1(SYNOPSYS_UNCONNECTED_110), .A2(
        \adder_sign/adder3/n81 ), .ZN(\adder_sign/adder3/n84 ) );
  XNOR2_X1 \adder_sign/adder3/U48  ( .A(n597), .B(1'b0), .ZN(
        \adder_sign/adder3/n83 ) );
  OAI22_X1 \adder_sign/adder3/U47  ( .A1(\adder_sign/adder3/n103 ), .A2(
        \adder_sign/adder3/n84 ), .B1(\adder_sign/adder3/n83 ), .B2(
        \adder_sign/adder3/n63 ), .ZN(sign_fixed[18]) );
  NOR2_X1 \adder_sign/adder3/U46  ( .A1(1'b0), .A2(n598), .ZN(
        \adder_sign/adder3/n85 ) );
  NOR2_X1 \adder_sign/adder3/U45  ( .A1(1'b0), .A2(n596), .ZN(
        \adder_sign/adder3/n78 ) );
  NOR2_X1 \adder_sign/adder3/U44  ( .A1(1'b0), .A2(n601), .ZN(
        \adder_sign/adder3/n96 ) );
  OAI21_X1 \adder_sign/adder3/U43  ( .B1(SYNOPSYS_UNCONNECTED_105), .B2(
        \adder_sign/adder3/n99 ), .A(\adder_sign/adder3/n61 ), .ZN(
        \adder_sign/adder3/n100 ) );
  XNOR2_X1 \adder_sign/adder3/U42  ( .A(n602), .B(1'b0), .ZN(
        \adder_sign/adder3/n102 ) );
  OAI21_X1 \adder_sign/adder3/U41  ( .B1(\adder_sign/adder3/n102 ), .B2(
        \adder_sign/adder3/n61 ), .A(\adder_sign/adder3/n100 ), .ZN(
        sign_fixed[23]) );
  INV_X1 \adder_sign/adder3/U40  ( .A(\adder_sign/adder3/n71 ), .ZN(
        SYNOPSYS_UNCONNECTED_106) );
  INV_X1 \adder_sign/adder3/U39  ( .A(\adder_sign/adder3/n70 ), .ZN(
        SYNOPSYS_UNCONNECTED_109) );
  INV_X1 \adder_sign/adder3/U38  ( .A(\adder_sign/adder3/n69 ), .ZN(
        SYNOPSYS_UNCONNECTED_111) );
  INV_X1 \adder_sign/adder3/U37  ( .A(\adder_sign/adder3/n99 ), .ZN(
        SYNOPSYS_UNCONNECTED_73) );
  INV_X1 \adder_sign/adder3/U36  ( .A(\adder_sign/adder3/n88 ), .ZN(
        SYNOPSYS_UNCONNECTED_76) );
  INV_X1 \adder_sign/adder3/U35  ( .A(\adder_sign/adder3/n75 ), .ZN(
        SYNOPSYS_UNCONNECTED_80) );
  INV_X1 \adder_sign/adder3/U34  ( .A(\adder_sign/adder3/n92 ), .ZN(
        SYNOPSYS_UNCONNECTED_75) );
  INV_X1 \adder_sign/adder3/U33  ( .A(\adder_sign/adder3/n81 ), .ZN(
        SYNOPSYS_UNCONNECTED_78) );
  INV_X1 \adder_sign/adder3/U32  ( .A(\adder_sign/adder3/n78 ), .ZN(
        SYNOPSYS_UNCONNECTED_79) );
  INV_X1 \adder_sign/adder3/U31  ( .A(\adder_sign/adder3/n96 ), .ZN(
        SYNOPSYS_UNCONNECTED_74) );
  INV_X1 \adder_sign/adder3/U30  ( .A(\adder_sign/adder3/n85 ), .ZN(
        SYNOPSYS_UNCONNECTED_77) );
  NOR2_X1 \adder_sign/adder3/U29  ( .A1(SYNOPSYS_UNCONNECTED_106), .A2(
        \adder_sign/adder3/n96 ), .ZN(\adder_sign/adder3/n97 ) );
  XNOR2_X1 \adder_sign/adder3/U28  ( .A(\adder_sign/adder3/n98 ), .B(
        \adder_sign/adder3/n97 ), .ZN(sign_fixed[22]) );
  NAND4_X1 \adder_sign/adder3/U27  ( .A1(SYNOPSYS_UNCONNECTED_77), .A2(
        SYNOPSYS_UNCONNECTED_76), .A3(SYNOPSYS_UNCONNECTED_75), .A4(
        SYNOPSYS_UNCONNECTED_74), .ZN(\adder_sign/adder3/n74 ) );
  NAND4_X1 \adder_sign/adder3/U26  ( .A1(SYNOPSYS_UNCONNECTED_73), .A2(
        SYNOPSYS_UNCONNECTED_80), .A3(SYNOPSYS_UNCONNECTED_79), .A4(
        SYNOPSYS_UNCONNECTED_78), .ZN(\adder_sign/adder3/n73 ) );
  NOR2_X1 \adder_sign/adder3/U25  ( .A1(SYNOPSYS_UNCONNECTED_111), .A2(
        \adder_sign/adder3/n78 ), .ZN(\adder_sign/adder3/n79 ) );
  XNOR2_X1 \adder_sign/adder3/U24  ( .A(\adder_sign/adder3/n67 ), .B(
        \adder_sign/adder3/n79 ), .ZN(sign_fixed[17]) );
  NOR2_X1 \adder_sign/adder3/U23  ( .A1(SYNOPSYS_UNCONNECTED_109), .A2(
        \adder_sign/adder3/n85 ), .ZN(\adder_sign/adder3/n86 ) );
  XNOR2_X1 \adder_sign/adder3/U22  ( .A(\adder_sign/adder3/n68 ), .B(
        \adder_sign/adder3/n86 ), .ZN(sign_fixed[19]) );
  AOI21_X1 \adder_sign/adder3/U21  ( .B1(\adder_sign/adder3/n90 ), .B2(
        SYNOPSYS_UNCONNECTED_76), .A(SYNOPSYS_UNCONNECTED_108), .ZN(
        \adder_sign/adder3/n94 ) );
  AOI21_X1 \adder_sign/adder3/U20  ( .B1(SYNOPSYS_UNCONNECTED_80), .B2(
        \adder_sign/n16 ), .A(SYNOPSYS_UNCONNECTED_112), .ZN(
        \adder_sign/adder3/n80 ) );
  OAI21_X1 \adder_sign/adder3/U19  ( .B1(\adder_sign/adder3/n87 ), .B2(
        \adder_sign/adder3/n85 ), .A(\adder_sign/adder3/n70 ), .ZN(
        \adder_sign/adder3/n90 ) );
  XNOR2_X1 \adder_sign/adder3/U18  ( .A(\adder_sign/adder3/n72 ), .B(
        \adder_sign/adder3/n60 ), .ZN(\adder_sign/adder3/overflow ) );
  INV_X1 \adder_sign/adder3/U17  ( .A(\adder_sign/adder3/n62 ), .ZN(
        \adder_sign/adder3/n104 ) );
  NOR2_X1 \adder_sign/adder3/U16  ( .A1(\adder_sign/adder3/n74 ), .A2(
        \adder_sign/adder3/n73 ), .ZN(\adder_sign/p2 ) );
  AOI21_X1 \adder_sign/adder3/U15  ( .B1(\adder_sign/adder3/n82 ), .B2(
        SYNOPSYS_UNCONNECTED_78), .A(SYNOPSYS_UNCONNECTED_110), .ZN(
        \adder_sign/adder3/n87 ) );
  AOI21_X1 \adder_sign/adder3/U14  ( .B1(\adder_sign/adder3/n60 ), .B2(
        SYNOPSYS_UNCONNECTED_73), .A(SYNOPSYS_UNCONNECTED_105), .ZN(
        \adder_sign/adder3/n72 ) );
  AOI21_X1 \adder_sign/adder3/U13  ( .B1(\adder_sign/adder3/n63 ), .B2(
        SYNOPSYS_UNCONNECTED_78), .A(SYNOPSYS_UNCONNECTED_110), .ZN(
        \adder_sign/adder3/n68 ) );
  AOI21_X1 \adder_sign/adder3/U12  ( .B1(SYNOPSYS_UNCONNECTED_80), .B2(
        \adder_sign/n16 ), .A(SYNOPSYS_UNCONNECTED_112), .ZN(
        \adder_sign/adder3/n67 ) );
  OAI21_X1 \adder_sign/adder3/U11  ( .B1(\adder_sign/adder3/n80 ), .B2(
        \adder_sign/adder3/n78 ), .A(\adder_sign/adder3/n69 ), .ZN(
        \adder_sign/adder3/n82 ) );
  INV_X1 \adder_sign/adder3/U10  ( .A(\adder_sign/adder3/n66 ), .ZN(
        \adder_sign/adder3/n98 ) );
  INV_X1 \adder_sign/adder3/U9  ( .A(SYNOPSYS_UNCONNECTED_107), .ZN(
        \adder_sign/adder3/n65 ) );
  OAI21_X1 \adder_sign/adder3/U8  ( .B1(\adder_sign/adder3/n92 ), .B2(
        \adder_sign/adder3/n94 ), .A(\adder_sign/adder3/n65 ), .ZN(
        \adder_sign/adder3/n66 ) );
  INV_X1 \adder_sign/adder3/U7  ( .A(\adder_sign/adder3/n64 ), .ZN(
        \adder_sign/g2 ) );
  AOI21_X1 \adder_sign/adder3/U6  ( .B1(SYNOPSYS_UNCONNECTED_73), .B2(
        \adder_sign/adder3/n101 ), .A(SYNOPSYS_UNCONNECTED_105), .ZN(
        \adder_sign/adder3/n64 ) );
  OAI21_X1 \adder_sign/adder3/U5  ( .B1(\adder_sign/adder3/n98 ), .B2(
        \adder_sign/adder3/n96 ), .A(\adder_sign/adder3/n71 ), .ZN(
        \adder_sign/adder3/n101 ) );
  OAI21_X1 \adder_sign/adder3/U4  ( .B1(\adder_sign/adder3/n80 ), .B2(
        \adder_sign/adder3/n78 ), .A(\adder_sign/adder3/n69 ), .ZN(
        \adder_sign/adder3/n63 ) );
  CLKBUF_X1 \adder_sign/adder3/U3  ( .A(\adder_sign/adder3/n94 ), .Z(
        \adder_sign/adder3/n62 ) );
  OAI21_X1 \adder_sign/adder3/U2  ( .B1(\adder_sign/adder3/n98 ), .B2(
        \adder_sign/adder3/n96 ), .A(\adder_sign/adder3/n71 ), .ZN(
        \adder_sign/adder3/n61 ) );
  OAI21_X1 \adder_sign/adder3/U1  ( .B1(\adder_sign/adder3/n98 ), .B2(
        \adder_sign/adder3/n96 ), .A(\adder_sign/adder3/n71 ), .ZN(
        \adder_sign/adder3/n60 ) );
  AND2_X1 \adder_sign/adder4/U71  ( .A1(1'b0), .A2(n603), .ZN(
        SYNOPSYS_UNCONNECTED_104) );
  AND2_X1 \adder_sign/adder4/U70  ( .A1(1'b0), .A2(n607), .ZN(
        SYNOPSYS_UNCONNECTED_100) );
  AND2_X1 \adder_sign/adder4/U69  ( .A1(1'b0), .A2(n605), .ZN(
        SYNOPSYS_UNCONNECTED_102) );
  AND2_X1 \adder_sign/adder4/U68  ( .A1(1'b0), .A2(n608), .ZN(
        SYNOPSYS_UNCONNECTED_99) );
  AND2_X1 \adder_sign/adder4/U67  ( .A1(n610), .A2(1'b0), .ZN(
        SYNOPSYS_UNCONNECTED_97) );
  NAND2_X1 \adder_sign/adder4/U66  ( .A1(1'b0), .A2(n609), .ZN(
        \adder_sign/adder4/n71 ) );
  NAND2_X1 \adder_sign/adder4/U65  ( .A1(1'b0), .A2(n606), .ZN(
        \adder_sign/adder4/n70 ) );
  NAND2_X1 \adder_sign/adder4/U64  ( .A1(1'b0), .A2(n604), .ZN(
        \adder_sign/adder4/n69 ) );
  XNOR2_X1 \adder_sign/adder4/U63  ( .A(\adder_sign/adder4/n72 ), .B(
        \adder_sign/adder4/n65 ), .ZN(div_sign_ovf) );
  NOR2_X1 \adder_sign/adder4/U62  ( .A1(1'b0), .A2(n610), .ZN(
        \adder_sign/adder4/n98 ) );
  NOR2_X1 \adder_sign/adder4/U61  ( .A1(1'b0), .A2(n607), .ZN(
        \adder_sign/adder4/n88 ) );
  NOR2_X1 \adder_sign/adder4/U60  ( .A1(1'b0), .A2(n603), .ZN(
        \adder_sign/adder4/n75 ) );
  NOR2_X1 \adder_sign/adder4/U59  ( .A1(1'b0), .A2(n608), .ZN(
        \adder_sign/adder4/n92 ) );
  NOR2_X1 \adder_sign/adder4/U58  ( .A1(1'b0), .A2(n605), .ZN(
        \adder_sign/adder4/n81 ) );
  NOR2_X1 \adder_sign/adder4/U57  ( .A1(1'b0), .A2(n604), .ZN(
        \adder_sign/adder4/n78 ) );
  NOR2_X1 \adder_sign/adder4/U56  ( .A1(1'b0), .A2(n609), .ZN(
        \adder_sign/adder4/n96 ) );
  NOR2_X1 \adder_sign/adder4/U55  ( .A1(1'b0), .A2(n606), .ZN(
        \adder_sign/adder4/n85 ) );
  INV_X1 \adder_sign/adder4/U54  ( .A(\adder_sign/adder4/n66 ), .ZN(
        \adder_sign/adder4/n102 ) );
  NOR2_X1 \adder_sign/adder4/U53  ( .A1(SYNOPSYS_UNCONNECTED_102), .A2(
        \adder_sign/adder4/n81 ), .ZN(\adder_sign/adder4/n84 ) );
  XNOR2_X1 \adder_sign/adder4/U52  ( .A(n605), .B(1'b0), .ZN(
        \adder_sign/adder4/n83 ) );
  OAI22_X1 \adder_sign/adder4/U51  ( .A1(\adder_sign/adder4/n102 ), .A2(
        \adder_sign/adder4/n84 ), .B1(\adder_sign/adder4/n83 ), .B2(
        \adder_sign/adder4/n66 ), .ZN(sign_fixed[26]) );
  OAI21_X1 \adder_sign/adder4/U50  ( .B1(SYNOPSYS_UNCONNECTED_104), .B2(
        \adder_sign/adder4/n75 ), .A(\adder_sign/n17 ), .ZN(
        \adder_sign/adder4/n76 ) );
  XNOR2_X1 \adder_sign/adder4/U49  ( .A(n603), .B(1'b0), .ZN(
        \adder_sign/adder4/n77 ) );
  OAI21_X1 \adder_sign/adder4/U48  ( .B1(\adder_sign/n17 ), .B2(
        \adder_sign/adder4/n77 ), .A(\adder_sign/adder4/n76 ), .ZN(
        sign_fixed[24]) );
  OAI21_X1 \adder_sign/adder4/U47  ( .B1(SYNOPSYS_UNCONNECTED_100), .B2(
        \adder_sign/adder4/n88 ), .A(\adder_sign/adder4/n61 ), .ZN(
        \adder_sign/adder4/n89 ) );
  XNOR2_X1 \adder_sign/adder4/U46  ( .A(n607), .B(1'b0), .ZN(
        \adder_sign/adder4/n91 ) );
  OAI21_X1 \adder_sign/adder4/U45  ( .B1(\adder_sign/adder4/n91 ), .B2(
        \adder_sign/adder4/n61 ), .A(\adder_sign/adder4/n89 ), .ZN(
        sign_fixed[28]) );
  OAI21_X1 \adder_sign/adder4/U44  ( .B1(SYNOPSYS_UNCONNECTED_97), .B2(
        \adder_sign/adder4/n98 ), .A(\adder_sign/adder4/n100 ), .ZN(
        \adder_sign/adder4/n99 ) );
  XNOR2_X1 \adder_sign/adder4/U43  ( .A(n610), .B(1'b0), .ZN(
        \adder_sign/adder4/n101 ) );
  NOR2_X1 \adder_sign/adder4/U42  ( .A1(SYNOPSYS_UNCONNECTED_99), .A2(
        \adder_sign/adder4/n92 ), .ZN(\adder_sign/adder4/n93 ) );
  XNOR2_X1 \adder_sign/adder4/U41  ( .A(n608), .B(1'b0), .ZN(
        \adder_sign/adder4/n95 ) );
  OAI22_X1 \adder_sign/adder4/U40  ( .A1(\adder_sign/adder4/n95 ), .A2(
        \adder_sign/adder4/n103 ), .B1(\adder_sign/adder4/n94 ), .B2(
        \adder_sign/adder4/n93 ), .ZN(sign_fixed[29]) );
  INV_X1 \adder_sign/adder4/U39  ( .A(\adder_sign/adder4/n70 ), .ZN(
        SYNOPSYS_UNCONNECTED_101) );
  INV_X1 \adder_sign/adder4/U38  ( .A(\adder_sign/adder4/n71 ), .ZN(
        SYNOPSYS_UNCONNECTED_98) );
  INV_X1 \adder_sign/adder4/U37  ( .A(\adder_sign/adder4/n69 ), .ZN(
        SYNOPSYS_UNCONNECTED_103) );
  INV_X1 \adder_sign/adder4/U36  ( .A(\adder_sign/adder4/n98 ), .ZN(
        SYNOPSYS_UNCONNECTED_65) );
  INV_X1 \adder_sign/adder4/U35  ( .A(\adder_sign/adder4/n88 ), .ZN(
        SYNOPSYS_UNCONNECTED_68) );
  INV_X1 \adder_sign/adder4/U34  ( .A(\adder_sign/adder4/n75 ), .ZN(
        SYNOPSYS_UNCONNECTED_72) );
  INV_X1 \adder_sign/adder4/U33  ( .A(\adder_sign/adder4/n92 ), .ZN(
        SYNOPSYS_UNCONNECTED_67) );
  INV_X1 \adder_sign/adder4/U32  ( .A(\adder_sign/adder4/n81 ), .ZN(
        SYNOPSYS_UNCONNECTED_70) );
  INV_X1 \adder_sign/adder4/U31  ( .A(\adder_sign/adder4/n78 ), .ZN(
        SYNOPSYS_UNCONNECTED_71) );
  INV_X1 \adder_sign/adder4/U30  ( .A(\adder_sign/adder4/n96 ), .ZN(
        SYNOPSYS_UNCONNECTED_66) );
  INV_X1 \adder_sign/adder4/U29  ( .A(\adder_sign/adder4/n85 ), .ZN(
        SYNOPSYS_UNCONNECTED_69) );
  NAND4_X1 \adder_sign/adder4/U28  ( .A1(SYNOPSYS_UNCONNECTED_69), .A2(
        SYNOPSYS_UNCONNECTED_68), .A3(SYNOPSYS_UNCONNECTED_67), .A4(
        SYNOPSYS_UNCONNECTED_66), .ZN(\adder_sign/adder4/n74 ) );
  NAND4_X1 \adder_sign/adder4/U27  ( .A1(SYNOPSYS_UNCONNECTED_65), .A2(
        SYNOPSYS_UNCONNECTED_72), .A3(SYNOPSYS_UNCONNECTED_71), .A4(
        SYNOPSYS_UNCONNECTED_70), .ZN(\adder_sign/adder4/n73 ) );
  AOI21_X1 \adder_sign/adder4/U26  ( .B1(\adder_sign/adder4/n65 ), .B2(
        SYNOPSYS_UNCONNECTED_65), .A(SYNOPSYS_UNCONNECTED_97), .ZN(
        \adder_sign/adder4/n72 ) );
  NOR2_X1 \adder_sign/adder4/U25  ( .A1(SYNOPSYS_UNCONNECTED_103), .A2(
        \adder_sign/adder4/n78 ), .ZN(\adder_sign/adder4/n79 ) );
  XNOR2_X1 \adder_sign/adder4/U24  ( .A(\adder_sign/adder4/n68 ), .B(
        \adder_sign/adder4/n79 ), .ZN(sign_fixed[25]) );
  NOR2_X1 \adder_sign/adder4/U23  ( .A1(SYNOPSYS_UNCONNECTED_101), .A2(
        \adder_sign/adder4/n85 ), .ZN(\adder_sign/adder4/n86 ) );
  XNOR2_X1 \adder_sign/adder4/U22  ( .A(\adder_sign/adder4/n67 ), .B(
        \adder_sign/adder4/n86 ), .ZN(sign_fixed[27]) );
  NOR2_X1 \adder_sign/adder4/U21  ( .A1(SYNOPSYS_UNCONNECTED_98), .A2(
        \adder_sign/adder4/n96 ), .ZN(\adder_sign/adder4/n97 ) );
  XNOR2_X1 \adder_sign/adder4/U20  ( .A(\adder_sign/adder4/n62 ), .B(
        \adder_sign/adder4/n97 ), .ZN(sign_fixed[30]) );
  AOI21_X1 \adder_sign/adder4/U19  ( .B1(\adder_sign/adder4/n90 ), .B2(
        SYNOPSYS_UNCONNECTED_68), .A(SYNOPSYS_UNCONNECTED_100), .ZN(
        \adder_sign/adder4/n94 ) );
  AOI21_X1 \adder_sign/adder4/U18  ( .B1(SYNOPSYS_UNCONNECTED_72), .B2(
        \adder_sign/n17 ), .A(SYNOPSYS_UNCONNECTED_104), .ZN(
        \adder_sign/adder4/n80 ) );
  OAI21_X1 \adder_sign/adder4/U17  ( .B1(\adder_sign/adder4/n87 ), .B2(
        \adder_sign/adder4/n85 ), .A(\adder_sign/adder4/n70 ), .ZN(
        \adder_sign/adder4/n90 ) );
  OAI21_X1 \adder_sign/adder4/U16  ( .B1(\adder_sign/adder4/n80 ), .B2(
        \adder_sign/adder4/n78 ), .A(\adder_sign/adder4/n69 ), .ZN(
        \adder_sign/adder4/n82 ) );
  INV_X1 \adder_sign/adder4/U15  ( .A(\adder_sign/adder4/n72 ), .ZN(
        \adder_sign/adder4/gen ) );
  NOR2_X1 \adder_sign/adder4/U14  ( .A1(\adder_sign/adder4/n74 ), .A2(
        \adder_sign/adder4/n73 ), .ZN(\adder_sign/adder4/prop ) );
  INV_X1 \adder_sign/adder4/U13  ( .A(\adder_sign/adder4/n94 ), .ZN(
        \adder_sign/adder4/n103 ) );
  AOI21_X1 \adder_sign/adder4/U12  ( .B1(\adder_sign/adder4/n82 ), .B2(
        SYNOPSYS_UNCONNECTED_70), .A(SYNOPSYS_UNCONNECTED_102), .ZN(
        \adder_sign/adder4/n87 ) );
  AOI21_X1 \adder_sign/adder4/U11  ( .B1(SYNOPSYS_UNCONNECTED_72), .B2(
        \adder_sign/n17 ), .A(SYNOPSYS_UNCONNECTED_104), .ZN(
        \adder_sign/adder4/n68 ) );
  AOI21_X1 \adder_sign/adder4/U10  ( .B1(\adder_sign/adder4/n66 ), .B2(
        SYNOPSYS_UNCONNECTED_70), .A(SYNOPSYS_UNCONNECTED_102), .ZN(
        \adder_sign/adder4/n67 ) );
  OAI21_X1 \adder_sign/adder4/U9  ( .B1(\adder_sign/adder4/n80 ), .B2(
        \adder_sign/adder4/n78 ), .A(\adder_sign/adder4/n69 ), .ZN(
        \adder_sign/adder4/n66 ) );
  CLKBUF_X1 \adder_sign/adder4/U8  ( .A(\adder_sign/adder4/n100 ), .Z(
        \adder_sign/adder4/n65 ) );
  INV_X1 \adder_sign/adder4/U7  ( .A(SYNOPSYS_UNCONNECTED_99), .ZN(
        \adder_sign/adder4/n63 ) );
  OAI21_X1 \adder_sign/adder4/U6  ( .B1(\adder_sign/adder4/n92 ), .B2(
        \adder_sign/adder4/n94 ), .A(\adder_sign/adder4/n63 ), .ZN(
        \adder_sign/adder4/n64 ) );
  INV_X1 \adder_sign/adder4/U5  ( .A(\adder_sign/adder4/n64 ), .ZN(
        \adder_sign/adder4/n62 ) );
  OAI21_X1 \adder_sign/adder4/U4  ( .B1(\adder_sign/adder4/n62 ), .B2(
        \adder_sign/adder4/n96 ), .A(\adder_sign/adder4/n71 ), .ZN(
        \adder_sign/adder4/n100 ) );
  CLKBUF_X1 \adder_sign/adder4/U3  ( .A(\adder_sign/adder4/n90 ), .Z(
        \adder_sign/adder4/n61 ) );
  NAND2_X1 \adder_sign/adder4/U2  ( .A1(\adder_sign/adder4/n60 ), .A2(
        \adder_sign/adder4/n99 ), .ZN(sign_fixed[31]) );
  OR2_X1 \adder_sign/adder4/U1  ( .A1(\adder_sign/adder4/n100 ), .A2(
        \adder_sign/adder4/n101 ), .ZN(\adder_sign/adder4/n60 ) );
  BUF_X1 \product_reg/U7  ( .A(n365), .Z(\product_reg/n2 ) );
  BUF_X1 \product_reg/U6  ( .A(n365), .Z(\product_reg/n6 ) );
  BUF_X1 \product_reg/U5  ( .A(n365), .Z(\product_reg/n5 ) );
  BUF_X1 \product_reg/U4  ( .A(n365), .Z(\product_reg/n4 ) );
  BUF_X1 \product_reg/U3  ( .A(n365), .Z(\product_reg/n3 ) );
  CLKBUF_X1 \product_reg/U2  ( .A(product_in[32]), .Z(\product_reg/n1 ) );
  BUF_X1 \product_reg/U1  ( .A(n365), .Z(\product_reg/n7 ) );
  INV_X1 \product_reg/memory_0__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_0__dff/n7 ) );
  NAND2_X1 \product_reg/memory_0__dff/U3  ( .A1(\product_reg/n2 ), .A2(
        product_in[0]), .ZN(\product_reg/memory_0__dff/n6 ) );
  OAI21_X1 \product_reg/memory_0__dff/U2  ( .B1(\product_reg/n2 ), .B2(
        \product_reg/memory_0__dff/n5 ), .A(\product_reg/memory_0__dff/n6 ), 
        .ZN(\product_reg/memory_0__dff/n1 ) );
  DFFR_X1 \product_reg/memory_0__dff/q_reg  ( .D(
        \product_reg/memory_0__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_0__dff/n7 ), .Q(product_out[0]), .QN(
        \product_reg/memory_0__dff/n5 ) );
  INV_X1 \product_reg/memory_1__dff/U6  ( .A(1'b0), .ZN(
        \product_reg/memory_1__dff/n10 ) );
  NAND2_X1 \product_reg/memory_1__dff/U5  ( .A1(\product_reg/n2 ), .A2(
        product_in[1]), .ZN(\product_reg/memory_1__dff/n9 ) );
  OAI21_X1 \product_reg/memory_1__dff/U4  ( .B1(\product_reg/n2 ), .B2(
        \product_reg/memory_1__dff/n6 ), .A(\product_reg/memory_1__dff/n9 ), 
        .ZN(\product_reg/memory_1__dff/n1 ) );
  INV_X1 \product_reg/memory_1__dff/U3  ( .A(\product_reg/memory_1__dff/n5 ), 
        .ZN(\product_reg/memory_1__dff/n6 ) );
  INV_X1 \product_reg/memory_1__dff/U2  ( .A(\product_reg/memory_1__dff/n8 ), 
        .ZN(product_out[1]) );
  DFFR_X1 \product_reg/memory_1__dff/q_reg  ( .D(
        \product_reg/memory_1__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_1__dff/n10 ), .Q(\product_reg/memory_1__dff/n5 ), 
        .QN(\product_reg/memory_1__dff/n8 ) );
  OAI21_X1 \product_reg/memory_2__dff/U7  ( .B1(\product_reg/n2 ), .B2(
        \product_reg/memory_2__dff/n7 ), .A(\product_reg/memory_2__dff/n9 ), 
        .ZN(\product_reg/memory_2__dff/n1 ) );
  INV_X1 \product_reg/memory_2__dff/U6  ( .A(1'b0), .ZN(
        \product_reg/memory_2__dff/n10 ) );
  NAND2_X1 \product_reg/memory_2__dff/U5  ( .A1(\product_reg/n2 ), .A2(
        product_in[2]), .ZN(\product_reg/memory_2__dff/n9 ) );
  INV_X1 \product_reg/memory_2__dff/U2  ( .A(\product_reg/memory_2__dff/n1 ), 
        .ZN(\product_reg/memory_2__dff/n4 ) );
  SDFFR_X1 \product_reg/memory_2__dff/q_reg  ( .D(1'b1), .SI(1'b0), .SE(
        \product_reg/memory_2__dff/n4 ), .CK(clock), .RN(
        \product_reg/memory_2__dff/n10 ), .Q(product_out[2]), .QN(
        \product_reg/memory_2__dff/n7 ) );
  INV_X1 \product_reg/memory_3__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_3__dff/n7 ) );
  NAND2_X1 \product_reg/memory_3__dff/U3  ( .A1(\product_reg/n2 ), .A2(
        product_in[3]), .ZN(\product_reg/memory_3__dff/n6 ) );
  OAI21_X1 \product_reg/memory_3__dff/U2  ( .B1(\product_reg/n2 ), .B2(
        \product_reg/memory_3__dff/n5 ), .A(\product_reg/memory_3__dff/n6 ), 
        .ZN(\product_reg/memory_3__dff/n1 ) );
  DFFR_X1 \product_reg/memory_3__dff/q_reg  ( .D(
        \product_reg/memory_3__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_3__dff/n7 ), .Q(product_out[3]), .QN(
        \product_reg/memory_3__dff/n5 ) );
  INV_X1 \product_reg/memory_4__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_4__dff/n7 ) );
  NAND2_X1 \product_reg/memory_4__dff/U3  ( .A1(\product_reg/n2 ), .A2(
        product_in[4]), .ZN(\product_reg/memory_4__dff/n6 ) );
  OAI21_X1 \product_reg/memory_4__dff/U2  ( .B1(\product_reg/n2 ), .B2(
        \product_reg/memory_4__dff/n5 ), .A(\product_reg/memory_4__dff/n6 ), 
        .ZN(\product_reg/memory_4__dff/n1 ) );
  DFFR_X1 \product_reg/memory_4__dff/q_reg  ( .D(
        \product_reg/memory_4__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_4__dff/n7 ), .Q(product_out[4]), .QN(
        \product_reg/memory_4__dff/n5 ) );
  INV_X1 \product_reg/memory_5__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_5__dff/n7 ) );
  NAND2_X1 \product_reg/memory_5__dff/U3  ( .A1(\product_reg/n2 ), .A2(
        product_in[5]), .ZN(\product_reg/memory_5__dff/n6 ) );
  OAI21_X1 \product_reg/memory_5__dff/U2  ( .B1(\product_reg/n2 ), .B2(
        \product_reg/memory_5__dff/n5 ), .A(\product_reg/memory_5__dff/n6 ), 
        .ZN(\product_reg/memory_5__dff/n1 ) );
  DFFR_X1 \product_reg/memory_5__dff/q_reg  ( .D(
        \product_reg/memory_5__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_5__dff/n7 ), .Q(product_out[5]), .QN(
        \product_reg/memory_5__dff/n5 ) );
  INV_X1 \product_reg/memory_6__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_6__dff/n7 ) );
  NAND2_X1 \product_reg/memory_6__dff/U3  ( .A1(\product_reg/n2 ), .A2(
        product_in[6]), .ZN(\product_reg/memory_6__dff/n6 ) );
  OAI21_X1 \product_reg/memory_6__dff/U2  ( .B1(\product_reg/n2 ), .B2(
        \product_reg/memory_6__dff/n5 ), .A(\product_reg/memory_6__dff/n6 ), 
        .ZN(\product_reg/memory_6__dff/n1 ) );
  DFFR_X1 \product_reg/memory_6__dff/q_reg  ( .D(
        \product_reg/memory_6__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_6__dff/n7 ), .Q(product_out[6]), .QN(
        \product_reg/memory_6__dff/n5 ) );
  INV_X1 \product_reg/memory_7__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_7__dff/n7 ) );
  NAND2_X1 \product_reg/memory_7__dff/U3  ( .A1(\product_reg/n2 ), .A2(
        product_in[7]), .ZN(\product_reg/memory_7__dff/n6 ) );
  OAI21_X1 \product_reg/memory_7__dff/U2  ( .B1(\product_reg/n2 ), .B2(
        \product_reg/memory_7__dff/n5 ), .A(\product_reg/memory_7__dff/n6 ), 
        .ZN(\product_reg/memory_7__dff/n1 ) );
  DFFR_X1 \product_reg/memory_7__dff/q_reg  ( .D(
        \product_reg/memory_7__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_7__dff/n7 ), .Q(product_out[7]), .QN(
        \product_reg/memory_7__dff/n5 ) );
  INV_X1 \product_reg/memory_8__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_8__dff/n7 ) );
  NAND2_X1 \product_reg/memory_8__dff/U3  ( .A1(\product_reg/n2 ), .A2(
        product_in[8]), .ZN(\product_reg/memory_8__dff/n6 ) );
  OAI21_X1 \product_reg/memory_8__dff/U2  ( .B1(\product_reg/n2 ), .B2(
        \product_reg/memory_8__dff/n5 ), .A(\product_reg/memory_8__dff/n6 ), 
        .ZN(\product_reg/memory_8__dff/n1 ) );
  DFFR_X1 \product_reg/memory_8__dff/q_reg  ( .D(
        \product_reg/memory_8__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_8__dff/n7 ), .Q(product_out[8]), .QN(
        \product_reg/memory_8__dff/n5 ) );
  INV_X1 \product_reg/memory_9__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_9__dff/n7 ) );
  NAND2_X1 \product_reg/memory_9__dff/U3  ( .A1(\product_reg/n2 ), .A2(
        product_in[9]), .ZN(\product_reg/memory_9__dff/n6 ) );
  OAI21_X1 \product_reg/memory_9__dff/U2  ( .B1(\product_reg/n2 ), .B2(
        \product_reg/memory_9__dff/n5 ), .A(\product_reg/memory_9__dff/n6 ), 
        .ZN(\product_reg/memory_9__dff/n1 ) );
  DFFR_X1 \product_reg/memory_9__dff/q_reg  ( .D(
        \product_reg/memory_9__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_9__dff/n7 ), .Q(product_out[9]), .QN(
        \product_reg/memory_9__dff/n5 ) );
  INV_X1 \product_reg/memory_10__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_10__dff/n7 ) );
  NAND2_X1 \product_reg/memory_10__dff/U3  ( .A1(\product_reg/n2 ), .A2(
        product_in[10]), .ZN(\product_reg/memory_10__dff/n6 ) );
  OAI21_X1 \product_reg/memory_10__dff/U2  ( .B1(\product_reg/n2 ), .B2(
        \product_reg/memory_10__dff/n5 ), .A(\product_reg/memory_10__dff/n6 ), 
        .ZN(\product_reg/memory_10__dff/n1 ) );
  DFFR_X1 \product_reg/memory_10__dff/q_reg  ( .D(
        \product_reg/memory_10__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_10__dff/n7 ), .Q(product_out[10]), .QN(
        \product_reg/memory_10__dff/n5 ) );
  INV_X1 \product_reg/memory_11__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_11__dff/n7 ) );
  NAND2_X1 \product_reg/memory_11__dff/U3  ( .A1(\product_reg/n2 ), .A2(
        product_in[11]), .ZN(\product_reg/memory_11__dff/n6 ) );
  OAI21_X1 \product_reg/memory_11__dff/U2  ( .B1(\product_reg/n2 ), .B2(
        \product_reg/memory_11__dff/n5 ), .A(\product_reg/memory_11__dff/n6 ), 
        .ZN(\product_reg/memory_11__dff/n1 ) );
  DFFR_X1 \product_reg/memory_11__dff/q_reg  ( .D(
        \product_reg/memory_11__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_11__dff/n7 ), .Q(product_out[11]), .QN(
        \product_reg/memory_11__dff/n5 ) );
  INV_X1 \product_reg/memory_12__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_12__dff/n7 ) );
  NAND2_X1 \product_reg/memory_12__dff/U3  ( .A1(\product_reg/n3 ), .A2(
        product_in[12]), .ZN(\product_reg/memory_12__dff/n6 ) );
  OAI21_X1 \product_reg/memory_12__dff/U2  ( .B1(\product_reg/n3 ), .B2(
        \product_reg/memory_12__dff/n5 ), .A(\product_reg/memory_12__dff/n6 ), 
        .ZN(\product_reg/memory_12__dff/n1 ) );
  DFFR_X1 \product_reg/memory_12__dff/q_reg  ( .D(
        \product_reg/memory_12__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_12__dff/n7 ), .Q(product_out[12]), .QN(
        \product_reg/memory_12__dff/n5 ) );
  INV_X1 \product_reg/memory_13__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_13__dff/n7 ) );
  NAND2_X1 \product_reg/memory_13__dff/U3  ( .A1(\product_reg/n3 ), .A2(
        product_in[13]), .ZN(\product_reg/memory_13__dff/n6 ) );
  OAI21_X1 \product_reg/memory_13__dff/U2  ( .B1(\product_reg/n3 ), .B2(
        \product_reg/memory_13__dff/n5 ), .A(\product_reg/memory_13__dff/n6 ), 
        .ZN(\product_reg/memory_13__dff/n1 ) );
  DFFR_X1 \product_reg/memory_13__dff/q_reg  ( .D(
        \product_reg/memory_13__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_13__dff/n7 ), .Q(product_out[13]), .QN(
        \product_reg/memory_13__dff/n5 ) );
  INV_X1 \product_reg/memory_14__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_14__dff/n7 ) );
  NAND2_X1 \product_reg/memory_14__dff/U3  ( .A1(\product_reg/n3 ), .A2(
        product_in[14]), .ZN(\product_reg/memory_14__dff/n6 ) );
  OAI21_X1 \product_reg/memory_14__dff/U2  ( .B1(\product_reg/n3 ), .B2(
        \product_reg/memory_14__dff/n5 ), .A(\product_reg/memory_14__dff/n6 ), 
        .ZN(\product_reg/memory_14__dff/n1 ) );
  DFFR_X1 \product_reg/memory_14__dff/q_reg  ( .D(
        \product_reg/memory_14__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_14__dff/n7 ), .Q(product_out[14]), .QN(
        \product_reg/memory_14__dff/n5 ) );
  INV_X1 \product_reg/memory_15__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_15__dff/n7 ) );
  NAND2_X1 \product_reg/memory_15__dff/U3  ( .A1(\product_reg/n3 ), .A2(
        product_in[15]), .ZN(\product_reg/memory_15__dff/n6 ) );
  OAI21_X1 \product_reg/memory_15__dff/U2  ( .B1(\product_reg/n3 ), .B2(
        \product_reg/memory_15__dff/n5 ), .A(\product_reg/memory_15__dff/n6 ), 
        .ZN(\product_reg/memory_15__dff/n1 ) );
  DFFR_X1 \product_reg/memory_15__dff/q_reg  ( .D(
        \product_reg/memory_15__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_15__dff/n7 ), .Q(product_out[15]), .QN(
        \product_reg/memory_15__dff/n5 ) );
  INV_X1 \product_reg/memory_16__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_16__dff/n7 ) );
  NAND2_X1 \product_reg/memory_16__dff/U3  ( .A1(\product_reg/n3 ), .A2(
        product_in[16]), .ZN(\product_reg/memory_16__dff/n6 ) );
  OAI21_X1 \product_reg/memory_16__dff/U2  ( .B1(\product_reg/n3 ), .B2(
        \product_reg/memory_16__dff/n5 ), .A(\product_reg/memory_16__dff/n6 ), 
        .ZN(\product_reg/memory_16__dff/n1 ) );
  DFFR_X1 \product_reg/memory_16__dff/q_reg  ( .D(
        \product_reg/memory_16__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_16__dff/n7 ), .Q(product_out[16]), .QN(
        \product_reg/memory_16__dff/n5 ) );
  INV_X1 \product_reg/memory_17__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_17__dff/n7 ) );
  NAND2_X1 \product_reg/memory_17__dff/U3  ( .A1(\product_reg/n3 ), .A2(
        product_in[17]), .ZN(\product_reg/memory_17__dff/n6 ) );
  OAI21_X1 \product_reg/memory_17__dff/U2  ( .B1(\product_reg/n3 ), .B2(
        \product_reg/memory_17__dff/n5 ), .A(\product_reg/memory_17__dff/n6 ), 
        .ZN(\product_reg/memory_17__dff/n1 ) );
  DFFR_X1 \product_reg/memory_17__dff/q_reg  ( .D(
        \product_reg/memory_17__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_17__dff/n7 ), .Q(product_out[17]), .QN(
        \product_reg/memory_17__dff/n5 ) );
  INV_X1 \product_reg/memory_18__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_18__dff/n7 ) );
  NAND2_X1 \product_reg/memory_18__dff/U3  ( .A1(\product_reg/n3 ), .A2(
        product_in[18]), .ZN(\product_reg/memory_18__dff/n6 ) );
  OAI21_X1 \product_reg/memory_18__dff/U2  ( .B1(\product_reg/n3 ), .B2(
        \product_reg/memory_18__dff/n5 ), .A(\product_reg/memory_18__dff/n6 ), 
        .ZN(\product_reg/memory_18__dff/n1 ) );
  DFFR_X1 \product_reg/memory_18__dff/q_reg  ( .D(
        \product_reg/memory_18__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_18__dff/n7 ), .Q(product_out[18]), .QN(
        \product_reg/memory_18__dff/n5 ) );
  INV_X1 \product_reg/memory_19__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_19__dff/n7 ) );
  NAND2_X1 \product_reg/memory_19__dff/U3  ( .A1(\product_reg/n3 ), .A2(
        product_in[19]), .ZN(\product_reg/memory_19__dff/n6 ) );
  OAI21_X1 \product_reg/memory_19__dff/U2  ( .B1(\product_reg/n3 ), .B2(
        \product_reg/memory_19__dff/n5 ), .A(\product_reg/memory_19__dff/n6 ), 
        .ZN(\product_reg/memory_19__dff/n1 ) );
  DFFR_X1 \product_reg/memory_19__dff/q_reg  ( .D(
        \product_reg/memory_19__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_19__dff/n7 ), .Q(product_out[19]), .QN(
        \product_reg/memory_19__dff/n5 ) );
  INV_X1 \product_reg/memory_20__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_20__dff/n7 ) );
  NAND2_X1 \product_reg/memory_20__dff/U3  ( .A1(\product_reg/n3 ), .A2(
        product_in[20]), .ZN(\product_reg/memory_20__dff/n6 ) );
  OAI21_X1 \product_reg/memory_20__dff/U2  ( .B1(\product_reg/n3 ), .B2(
        \product_reg/memory_20__dff/n5 ), .A(\product_reg/memory_20__dff/n6 ), 
        .ZN(\product_reg/memory_20__dff/n1 ) );
  DFFR_X1 \product_reg/memory_20__dff/q_reg  ( .D(
        \product_reg/memory_20__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_20__dff/n7 ), .Q(product_out[20]), .QN(
        \product_reg/memory_20__dff/n5 ) );
  INV_X1 \product_reg/memory_21__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_21__dff/n7 ) );
  NAND2_X1 \product_reg/memory_21__dff/U3  ( .A1(\product_reg/n3 ), .A2(
        product_in[21]), .ZN(\product_reg/memory_21__dff/n6 ) );
  OAI21_X1 \product_reg/memory_21__dff/U2  ( .B1(\product_reg/n3 ), .B2(
        \product_reg/memory_21__dff/n5 ), .A(\product_reg/memory_21__dff/n6 ), 
        .ZN(\product_reg/memory_21__dff/n1 ) );
  DFFR_X1 \product_reg/memory_21__dff/q_reg  ( .D(
        \product_reg/memory_21__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_21__dff/n7 ), .Q(product_out[21]), .QN(
        \product_reg/memory_21__dff/n5 ) );
  INV_X1 \product_reg/memory_22__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_22__dff/n7 ) );
  NAND2_X1 \product_reg/memory_22__dff/U3  ( .A1(\product_reg/n3 ), .A2(
        product_in[22]), .ZN(\product_reg/memory_22__dff/n6 ) );
  OAI21_X1 \product_reg/memory_22__dff/U2  ( .B1(\product_reg/n3 ), .B2(
        \product_reg/memory_22__dff/n5 ), .A(\product_reg/memory_22__dff/n6 ), 
        .ZN(\product_reg/memory_22__dff/n1 ) );
  DFFR_X1 \product_reg/memory_22__dff/q_reg  ( .D(
        \product_reg/memory_22__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_22__dff/n7 ), .Q(product_out[22]), .QN(
        \product_reg/memory_22__dff/n5 ) );
  INV_X1 \product_reg/memory_23__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_23__dff/n7 ) );
  NAND2_X1 \product_reg/memory_23__dff/U3  ( .A1(\product_reg/n3 ), .A2(
        product_in[23]), .ZN(\product_reg/memory_23__dff/n6 ) );
  OAI21_X1 \product_reg/memory_23__dff/U2  ( .B1(\product_reg/n3 ), .B2(
        \product_reg/memory_23__dff/n5 ), .A(\product_reg/memory_23__dff/n6 ), 
        .ZN(\product_reg/memory_23__dff/n1 ) );
  DFFR_X1 \product_reg/memory_23__dff/q_reg  ( .D(
        \product_reg/memory_23__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_23__dff/n7 ), .Q(product_out[23]), .QN(
        \product_reg/memory_23__dff/n5 ) );
  INV_X1 \product_reg/memory_24__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_24__dff/n7 ) );
  NAND2_X1 \product_reg/memory_24__dff/U3  ( .A1(\product_reg/n4 ), .A2(
        product_in[24]), .ZN(\product_reg/memory_24__dff/n6 ) );
  OAI21_X1 \product_reg/memory_24__dff/U2  ( .B1(\product_reg/n4 ), .B2(
        \product_reg/memory_24__dff/n5 ), .A(\product_reg/memory_24__dff/n6 ), 
        .ZN(\product_reg/memory_24__dff/n1 ) );
  DFFR_X1 \product_reg/memory_24__dff/q_reg  ( .D(
        \product_reg/memory_24__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_24__dff/n7 ), .Q(product_out[24]), .QN(
        \product_reg/memory_24__dff/n5 ) );
  INV_X1 \product_reg/memory_25__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_25__dff/n7 ) );
  NAND2_X1 \product_reg/memory_25__dff/U3  ( .A1(\product_reg/n4 ), .A2(
        product_in[25]), .ZN(\product_reg/memory_25__dff/n6 ) );
  OAI21_X1 \product_reg/memory_25__dff/U2  ( .B1(\product_reg/n4 ), .B2(
        \product_reg/memory_25__dff/n5 ), .A(\product_reg/memory_25__dff/n6 ), 
        .ZN(\product_reg/memory_25__dff/n1 ) );
  DFFR_X1 \product_reg/memory_25__dff/q_reg  ( .D(
        \product_reg/memory_25__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_25__dff/n7 ), .Q(product_out[25]), .QN(
        \product_reg/memory_25__dff/n5 ) );
  INV_X1 \product_reg/memory_26__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_26__dff/n7 ) );
  NAND2_X1 \product_reg/memory_26__dff/U3  ( .A1(\product_reg/n4 ), .A2(
        product_in[26]), .ZN(\product_reg/memory_26__dff/n6 ) );
  OAI21_X1 \product_reg/memory_26__dff/U2  ( .B1(\product_reg/n4 ), .B2(
        \product_reg/memory_26__dff/n5 ), .A(\product_reg/memory_26__dff/n6 ), 
        .ZN(\product_reg/memory_26__dff/n1 ) );
  DFFR_X1 \product_reg/memory_26__dff/q_reg  ( .D(
        \product_reg/memory_26__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_26__dff/n7 ), .Q(product_out[26]), .QN(
        \product_reg/memory_26__dff/n5 ) );
  INV_X1 \product_reg/memory_27__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_27__dff/n7 ) );
  NAND2_X1 \product_reg/memory_27__dff/U3  ( .A1(\product_reg/n4 ), .A2(
        product_in[27]), .ZN(\product_reg/memory_27__dff/n6 ) );
  OAI21_X1 \product_reg/memory_27__dff/U2  ( .B1(\product_reg/n4 ), .B2(
        \product_reg/memory_27__dff/n5 ), .A(\product_reg/memory_27__dff/n6 ), 
        .ZN(\product_reg/memory_27__dff/n1 ) );
  DFFR_X1 \product_reg/memory_27__dff/q_reg  ( .D(
        \product_reg/memory_27__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_27__dff/n7 ), .Q(product_out[27]), .QN(
        \product_reg/memory_27__dff/n5 ) );
  INV_X1 \product_reg/memory_28__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_28__dff/n7 ) );
  NAND2_X1 \product_reg/memory_28__dff/U3  ( .A1(\product_reg/n4 ), .A2(
        product_in[28]), .ZN(\product_reg/memory_28__dff/n6 ) );
  OAI21_X1 \product_reg/memory_28__dff/U2  ( .B1(\product_reg/n4 ), .B2(
        \product_reg/memory_28__dff/n5 ), .A(\product_reg/memory_28__dff/n6 ), 
        .ZN(\product_reg/memory_28__dff/n1 ) );
  DFFR_X1 \product_reg/memory_28__dff/q_reg  ( .D(
        \product_reg/memory_28__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_28__dff/n7 ), .Q(product_out[28]), .QN(
        \product_reg/memory_28__dff/n5 ) );
  INV_X1 \product_reg/memory_29__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_29__dff/n7 ) );
  NAND2_X1 \product_reg/memory_29__dff/U3  ( .A1(\product_reg/n4 ), .A2(
        product_in[29]), .ZN(\product_reg/memory_29__dff/n6 ) );
  OAI21_X1 \product_reg/memory_29__dff/U2  ( .B1(\product_reg/n4 ), .B2(
        \product_reg/memory_29__dff/n5 ), .A(\product_reg/memory_29__dff/n6 ), 
        .ZN(\product_reg/memory_29__dff/n1 ) );
  DFFR_X1 \product_reg/memory_29__dff/q_reg  ( .D(
        \product_reg/memory_29__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_29__dff/n7 ), .Q(product_out[29]), .QN(
        \product_reg/memory_29__dff/n5 ) );
  INV_X1 \product_reg/memory_30__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_30__dff/n7 ) );
  NAND2_X1 \product_reg/memory_30__dff/U3  ( .A1(\product_reg/n4 ), .A2(
        product_in[30]), .ZN(\product_reg/memory_30__dff/n6 ) );
  OAI21_X1 \product_reg/memory_30__dff/U2  ( .B1(\product_reg/n4 ), .B2(
        \product_reg/memory_30__dff/n5 ), .A(\product_reg/memory_30__dff/n6 ), 
        .ZN(\product_reg/memory_30__dff/n1 ) );
  DFFR_X1 \product_reg/memory_30__dff/q_reg  ( .D(
        \product_reg/memory_30__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_30__dff/n7 ), .Q(product_out[30]), .QN(
        \product_reg/memory_30__dff/n5 ) );
  INV_X1 \product_reg/memory_31__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_31__dff/n7 ) );
  NAND2_X1 \product_reg/memory_31__dff/U3  ( .A1(\product_reg/n4 ), .A2(
        product_in[31]), .ZN(\product_reg/memory_31__dff/n6 ) );
  OAI21_X1 \product_reg/memory_31__dff/U2  ( .B1(\product_reg/n4 ), .B2(
        \product_reg/memory_31__dff/n5 ), .A(\product_reg/memory_31__dff/n6 ), 
        .ZN(\product_reg/memory_31__dff/n1 ) );
  DFFR_X1 \product_reg/memory_31__dff/q_reg  ( .D(
        \product_reg/memory_31__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_31__dff/n7 ), .Q(product_out[31]), .QN(
        \product_reg/memory_31__dff/n5 ) );
  INV_X1 \product_reg/memory_32__dff/U3  ( .A(1'b0), .ZN(
        \product_reg/memory_32__dff/n3 ) );
  MUX2_X1 \product_reg/memory_32__dff/U2  ( .A(product_out[32]), .B(
        \product_reg/n1 ), .S(\product_reg/n4 ), .Z(
        \product_reg/memory_32__dff/n1 ) );
  DFFR_X1 \product_reg/memory_32__dff/q_reg  ( .D(
        \product_reg/memory_32__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_32__dff/n3 ), .Q(product_out[32]), .QN() );
  INV_X1 \product_reg/memory_33__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_33__dff/n7 ) );
  NAND2_X1 \product_reg/memory_33__dff/U3  ( .A1(\product_reg/n4 ), .A2(
        product_in[33]), .ZN(\product_reg/memory_33__dff/n6 ) );
  OAI21_X1 \product_reg/memory_33__dff/U2  ( .B1(\product_reg/n4 ), .B2(
        \product_reg/memory_33__dff/n5 ), .A(\product_reg/memory_33__dff/n6 ), 
        .ZN(\product_reg/memory_33__dff/n1 ) );
  DFFR_X1 \product_reg/memory_33__dff/q_reg  ( .D(
        \product_reg/memory_33__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_33__dff/n7 ), .Q(product_out[33]), .QN(
        \product_reg/memory_33__dff/n5 ) );
  INV_X1 \product_reg/memory_34__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_34__dff/n7 ) );
  NAND2_X1 \product_reg/memory_34__dff/U3  ( .A1(\product_reg/n4 ), .A2(
        product_in[34]), .ZN(\product_reg/memory_34__dff/n6 ) );
  OAI21_X1 \product_reg/memory_34__dff/U2  ( .B1(\product_reg/n4 ), .B2(
        \product_reg/memory_34__dff/n5 ), .A(\product_reg/memory_34__dff/n6 ), 
        .ZN(\product_reg/memory_34__dff/n1 ) );
  DFFR_X1 \product_reg/memory_34__dff/q_reg  ( .D(
        \product_reg/memory_34__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_34__dff/n7 ), .Q(product_out[34]), .QN(
        \product_reg/memory_34__dff/n5 ) );
  INV_X1 \product_reg/memory_35__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_35__dff/n7 ) );
  NAND2_X1 \product_reg/memory_35__dff/U3  ( .A1(\product_reg/n4 ), .A2(
        product_in[35]), .ZN(\product_reg/memory_35__dff/n6 ) );
  OAI21_X1 \product_reg/memory_35__dff/U2  ( .B1(\product_reg/n4 ), .B2(
        \product_reg/memory_35__dff/n5 ), .A(\product_reg/memory_35__dff/n6 ), 
        .ZN(\product_reg/memory_35__dff/n1 ) );
  DFFR_X1 \product_reg/memory_35__dff/q_reg  ( .D(
        \product_reg/memory_35__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_35__dff/n7 ), .Q(product_out[35]), .QN(
        \product_reg/memory_35__dff/n5 ) );
  INV_X1 \product_reg/memory_36__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_36__dff/n7 ) );
  NAND2_X1 \product_reg/memory_36__dff/U3  ( .A1(\product_reg/n5 ), .A2(
        product_in[36]), .ZN(\product_reg/memory_36__dff/n6 ) );
  OAI21_X1 \product_reg/memory_36__dff/U2  ( .B1(\product_reg/n5 ), .B2(
        \product_reg/memory_36__dff/n5 ), .A(\product_reg/memory_36__dff/n6 ), 
        .ZN(\product_reg/memory_36__dff/n1 ) );
  DFFR_X1 \product_reg/memory_36__dff/q_reg  ( .D(
        \product_reg/memory_36__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_36__dff/n7 ), .Q(product_out[36]), .QN(
        \product_reg/memory_36__dff/n5 ) );
  INV_X1 \product_reg/memory_37__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_37__dff/n7 ) );
  NAND2_X1 \product_reg/memory_37__dff/U3  ( .A1(\product_reg/n5 ), .A2(
        product_in[37]), .ZN(\product_reg/memory_37__dff/n6 ) );
  OAI21_X1 \product_reg/memory_37__dff/U2  ( .B1(\product_reg/n5 ), .B2(
        \product_reg/memory_37__dff/n5 ), .A(\product_reg/memory_37__dff/n6 ), 
        .ZN(\product_reg/memory_37__dff/n1 ) );
  DFFR_X1 \product_reg/memory_37__dff/q_reg  ( .D(
        \product_reg/memory_37__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_37__dff/n7 ), .Q(product_out[37]), .QN(
        \product_reg/memory_37__dff/n5 ) );
  INV_X1 \product_reg/memory_38__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_38__dff/n7 ) );
  NAND2_X1 \product_reg/memory_38__dff/U3  ( .A1(\product_reg/n5 ), .A2(
        product_in[38]), .ZN(\product_reg/memory_38__dff/n6 ) );
  OAI21_X1 \product_reg/memory_38__dff/U2  ( .B1(\product_reg/n5 ), .B2(
        \product_reg/memory_38__dff/n5 ), .A(\product_reg/memory_38__dff/n6 ), 
        .ZN(\product_reg/memory_38__dff/n1 ) );
  DFFR_X1 \product_reg/memory_38__dff/q_reg  ( .D(
        \product_reg/memory_38__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_38__dff/n7 ), .Q(product_out[38]), .QN(
        \product_reg/memory_38__dff/n5 ) );
  INV_X1 \product_reg/memory_39__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_39__dff/n7 ) );
  NAND2_X1 \product_reg/memory_39__dff/U3  ( .A1(\product_reg/n5 ), .A2(
        product_in[39]), .ZN(\product_reg/memory_39__dff/n6 ) );
  OAI21_X1 \product_reg/memory_39__dff/U2  ( .B1(\product_reg/n5 ), .B2(
        \product_reg/memory_39__dff/n5 ), .A(\product_reg/memory_39__dff/n6 ), 
        .ZN(\product_reg/memory_39__dff/n1 ) );
  DFFR_X1 \product_reg/memory_39__dff/q_reg  ( .D(
        \product_reg/memory_39__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_39__dff/n7 ), .Q(product_out[39]), .QN(
        \product_reg/memory_39__dff/n5 ) );
  INV_X1 \product_reg/memory_40__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_40__dff/n7 ) );
  NAND2_X1 \product_reg/memory_40__dff/U3  ( .A1(\product_reg/n5 ), .A2(
        product_in[40]), .ZN(\product_reg/memory_40__dff/n6 ) );
  OAI21_X1 \product_reg/memory_40__dff/U2  ( .B1(\product_reg/n5 ), .B2(
        \product_reg/memory_40__dff/n5 ), .A(\product_reg/memory_40__dff/n6 ), 
        .ZN(\product_reg/memory_40__dff/n1 ) );
  DFFR_X1 \product_reg/memory_40__dff/q_reg  ( .D(
        \product_reg/memory_40__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_40__dff/n7 ), .Q(product_out[40]), .QN(
        \product_reg/memory_40__dff/n5 ) );
  INV_X1 \product_reg/memory_41__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_41__dff/n7 ) );
  NAND2_X1 \product_reg/memory_41__dff/U3  ( .A1(\product_reg/n5 ), .A2(
        product_in[41]), .ZN(\product_reg/memory_41__dff/n6 ) );
  OAI21_X1 \product_reg/memory_41__dff/U2  ( .B1(\product_reg/n5 ), .B2(
        \product_reg/memory_41__dff/n5 ), .A(\product_reg/memory_41__dff/n6 ), 
        .ZN(\product_reg/memory_41__dff/n1 ) );
  DFFR_X1 \product_reg/memory_41__dff/q_reg  ( .D(
        \product_reg/memory_41__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_41__dff/n7 ), .Q(product_out[41]), .QN(
        \product_reg/memory_41__dff/n5 ) );
  INV_X1 \product_reg/memory_42__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_42__dff/n7 ) );
  NAND2_X1 \product_reg/memory_42__dff/U3  ( .A1(\product_reg/n5 ), .A2(
        product_in[42]), .ZN(\product_reg/memory_42__dff/n6 ) );
  OAI21_X1 \product_reg/memory_42__dff/U2  ( .B1(\product_reg/n5 ), .B2(
        \product_reg/memory_42__dff/n5 ), .A(\product_reg/memory_42__dff/n6 ), 
        .ZN(\product_reg/memory_42__dff/n1 ) );
  DFFR_X1 \product_reg/memory_42__dff/q_reg  ( .D(
        \product_reg/memory_42__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_42__dff/n7 ), .Q(product_out[42]), .QN(
        \product_reg/memory_42__dff/n5 ) );
  INV_X1 \product_reg/memory_43__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_43__dff/n7 ) );
  NAND2_X1 \product_reg/memory_43__dff/U3  ( .A1(\product_reg/n5 ), .A2(
        product_in[43]), .ZN(\product_reg/memory_43__dff/n6 ) );
  OAI21_X1 \product_reg/memory_43__dff/U2  ( .B1(\product_reg/n5 ), .B2(
        \product_reg/memory_43__dff/n5 ), .A(\product_reg/memory_43__dff/n6 ), 
        .ZN(\product_reg/memory_43__dff/n1 ) );
  DFFR_X1 \product_reg/memory_43__dff/q_reg  ( .D(
        \product_reg/memory_43__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_43__dff/n7 ), .Q(product_out[43]), .QN(
        \product_reg/memory_43__dff/n5 ) );
  INV_X1 \product_reg/memory_44__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_44__dff/n7 ) );
  NAND2_X1 \product_reg/memory_44__dff/U3  ( .A1(\product_reg/n5 ), .A2(
        product_in[44]), .ZN(\product_reg/memory_44__dff/n6 ) );
  OAI21_X1 \product_reg/memory_44__dff/U2  ( .B1(\product_reg/n5 ), .B2(
        \product_reg/memory_44__dff/n5 ), .A(\product_reg/memory_44__dff/n6 ), 
        .ZN(\product_reg/memory_44__dff/n1 ) );
  DFFR_X1 \product_reg/memory_44__dff/q_reg  ( .D(
        \product_reg/memory_44__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_44__dff/n7 ), .Q(product_out[44]), .QN(
        \product_reg/memory_44__dff/n5 ) );
  INV_X1 \product_reg/memory_45__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_45__dff/n7 ) );
  NAND2_X1 \product_reg/memory_45__dff/U3  ( .A1(\product_reg/n5 ), .A2(
        product_in[45]), .ZN(\product_reg/memory_45__dff/n6 ) );
  OAI21_X1 \product_reg/memory_45__dff/U2  ( .B1(\product_reg/n5 ), .B2(
        \product_reg/memory_45__dff/n5 ), .A(\product_reg/memory_45__dff/n6 ), 
        .ZN(\product_reg/memory_45__dff/n1 ) );
  DFFR_X1 \product_reg/memory_45__dff/q_reg  ( .D(
        \product_reg/memory_45__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_45__dff/n7 ), .Q(product_out[45]), .QN(
        \product_reg/memory_45__dff/n5 ) );
  INV_X1 \product_reg/memory_46__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_46__dff/n7 ) );
  NAND2_X1 \product_reg/memory_46__dff/U3  ( .A1(\product_reg/n5 ), .A2(
        product_in[46]), .ZN(\product_reg/memory_46__dff/n6 ) );
  OAI21_X1 \product_reg/memory_46__dff/U2  ( .B1(\product_reg/n5 ), .B2(
        \product_reg/memory_46__dff/n5 ), .A(\product_reg/memory_46__dff/n6 ), 
        .ZN(\product_reg/memory_46__dff/n1 ) );
  DFFR_X1 \product_reg/memory_46__dff/q_reg  ( .D(
        \product_reg/memory_46__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_46__dff/n7 ), .Q(product_out[46]), .QN(
        \product_reg/memory_46__dff/n5 ) );
  INV_X1 \product_reg/memory_47__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_47__dff/n7 ) );
  NAND2_X1 \product_reg/memory_47__dff/U3  ( .A1(\product_reg/n5 ), .A2(
        product_in[47]), .ZN(\product_reg/memory_47__dff/n6 ) );
  OAI21_X1 \product_reg/memory_47__dff/U2  ( .B1(\product_reg/n5 ), .B2(
        \product_reg/memory_47__dff/n5 ), .A(\product_reg/memory_47__dff/n6 ), 
        .ZN(\product_reg/memory_47__dff/n1 ) );
  DFFR_X1 \product_reg/memory_47__dff/q_reg  ( .D(
        \product_reg/memory_47__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_47__dff/n7 ), .Q(product_out[47]), .QN(
        \product_reg/memory_47__dff/n5 ) );
  INV_X1 \product_reg/memory_48__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_48__dff/n7 ) );
  NAND2_X1 \product_reg/memory_48__dff/U3  ( .A1(\product_reg/n6 ), .A2(
        product_in[48]), .ZN(\product_reg/memory_48__dff/n6 ) );
  OAI21_X1 \product_reg/memory_48__dff/U2  ( .B1(\product_reg/n6 ), .B2(
        \product_reg/memory_48__dff/n5 ), .A(\product_reg/memory_48__dff/n6 ), 
        .ZN(\product_reg/memory_48__dff/n1 ) );
  DFFR_X1 \product_reg/memory_48__dff/q_reg  ( .D(
        \product_reg/memory_48__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_48__dff/n7 ), .Q(product_out[48]), .QN(
        \product_reg/memory_48__dff/n5 ) );
  INV_X1 \product_reg/memory_49__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_49__dff/n7 ) );
  NAND2_X1 \product_reg/memory_49__dff/U3  ( .A1(\product_reg/n6 ), .A2(
        product_in[49]), .ZN(\product_reg/memory_49__dff/n6 ) );
  OAI21_X1 \product_reg/memory_49__dff/U2  ( .B1(\product_reg/n6 ), .B2(
        \product_reg/memory_49__dff/n5 ), .A(\product_reg/memory_49__dff/n6 ), 
        .ZN(\product_reg/memory_49__dff/n1 ) );
  DFFR_X1 \product_reg/memory_49__dff/q_reg  ( .D(
        \product_reg/memory_49__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_49__dff/n7 ), .Q(product_out[49]), .QN(
        \product_reg/memory_49__dff/n5 ) );
  INV_X1 \product_reg/memory_50__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_50__dff/n7 ) );
  NAND2_X1 \product_reg/memory_50__dff/U3  ( .A1(\product_reg/n6 ), .A2(
        product_in[50]), .ZN(\product_reg/memory_50__dff/n6 ) );
  OAI21_X1 \product_reg/memory_50__dff/U2  ( .B1(\product_reg/n6 ), .B2(
        \product_reg/memory_50__dff/n5 ), .A(\product_reg/memory_50__dff/n6 ), 
        .ZN(\product_reg/memory_50__dff/n1 ) );
  DFFR_X1 \product_reg/memory_50__dff/q_reg  ( .D(
        \product_reg/memory_50__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_50__dff/n7 ), .Q(product_out[50]), .QN(
        \product_reg/memory_50__dff/n5 ) );
  INV_X1 \product_reg/memory_51__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_51__dff/n7 ) );
  NAND2_X1 \product_reg/memory_51__dff/U3  ( .A1(\product_reg/n6 ), .A2(
        product_in[51]), .ZN(\product_reg/memory_51__dff/n6 ) );
  OAI21_X1 \product_reg/memory_51__dff/U2  ( .B1(\product_reg/n6 ), .B2(
        \product_reg/memory_51__dff/n5 ), .A(\product_reg/memory_51__dff/n6 ), 
        .ZN(\product_reg/memory_51__dff/n1 ) );
  DFFR_X1 \product_reg/memory_51__dff/q_reg  ( .D(
        \product_reg/memory_51__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_51__dff/n7 ), .Q(product_out[51]), .QN(
        \product_reg/memory_51__dff/n5 ) );
  INV_X1 \product_reg/memory_52__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_52__dff/n7 ) );
  NAND2_X1 \product_reg/memory_52__dff/U3  ( .A1(\product_reg/n6 ), .A2(
        product_in[52]), .ZN(\product_reg/memory_52__dff/n6 ) );
  OAI21_X1 \product_reg/memory_52__dff/U2  ( .B1(\product_reg/n6 ), .B2(
        \product_reg/memory_52__dff/n5 ), .A(\product_reg/memory_52__dff/n6 ), 
        .ZN(\product_reg/memory_52__dff/n1 ) );
  DFFR_X1 \product_reg/memory_52__dff/q_reg  ( .D(
        \product_reg/memory_52__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_52__dff/n7 ), .Q(product_out[52]), .QN(
        \product_reg/memory_52__dff/n5 ) );
  INV_X1 \product_reg/memory_53__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_53__dff/n7 ) );
  NAND2_X1 \product_reg/memory_53__dff/U3  ( .A1(\product_reg/n6 ), .A2(
        product_in[53]), .ZN(\product_reg/memory_53__dff/n6 ) );
  OAI21_X1 \product_reg/memory_53__dff/U2  ( .B1(\product_reg/n6 ), .B2(
        \product_reg/memory_53__dff/n5 ), .A(\product_reg/memory_53__dff/n6 ), 
        .ZN(\product_reg/memory_53__dff/n1 ) );
  DFFR_X1 \product_reg/memory_53__dff/q_reg  ( .D(
        \product_reg/memory_53__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_53__dff/n7 ), .Q(product_out[53]), .QN(
        \product_reg/memory_53__dff/n5 ) );
  INV_X1 \product_reg/memory_54__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_54__dff/n7 ) );
  NAND2_X1 \product_reg/memory_54__dff/U3  ( .A1(\product_reg/n6 ), .A2(
        product_in[54]), .ZN(\product_reg/memory_54__dff/n6 ) );
  OAI21_X1 \product_reg/memory_54__dff/U2  ( .B1(\product_reg/n6 ), .B2(
        \product_reg/memory_54__dff/n5 ), .A(\product_reg/memory_54__dff/n6 ), 
        .ZN(\product_reg/memory_54__dff/n1 ) );
  DFFR_X1 \product_reg/memory_54__dff/q_reg  ( .D(
        \product_reg/memory_54__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_54__dff/n7 ), .Q(product_out[54]), .QN(
        \product_reg/memory_54__dff/n5 ) );
  INV_X1 \product_reg/memory_55__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_55__dff/n7 ) );
  NAND2_X1 \product_reg/memory_55__dff/U3  ( .A1(\product_reg/n6 ), .A2(
        product_in[55]), .ZN(\product_reg/memory_55__dff/n6 ) );
  OAI21_X1 \product_reg/memory_55__dff/U2  ( .B1(\product_reg/n6 ), .B2(
        \product_reg/memory_55__dff/n5 ), .A(\product_reg/memory_55__dff/n6 ), 
        .ZN(\product_reg/memory_55__dff/n1 ) );
  DFFR_X1 \product_reg/memory_55__dff/q_reg  ( .D(
        \product_reg/memory_55__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_55__dff/n7 ), .Q(product_out[55]), .QN(
        \product_reg/memory_55__dff/n5 ) );
  INV_X1 \product_reg/memory_56__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_56__dff/n7 ) );
  NAND2_X1 \product_reg/memory_56__dff/U3  ( .A1(\product_reg/n6 ), .A2(
        product_in[56]), .ZN(\product_reg/memory_56__dff/n6 ) );
  OAI21_X1 \product_reg/memory_56__dff/U2  ( .B1(\product_reg/n6 ), .B2(
        \product_reg/memory_56__dff/n5 ), .A(\product_reg/memory_56__dff/n6 ), 
        .ZN(\product_reg/memory_56__dff/n1 ) );
  DFFR_X1 \product_reg/memory_56__dff/q_reg  ( .D(
        \product_reg/memory_56__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_56__dff/n7 ), .Q(product_out[56]), .QN(
        \product_reg/memory_56__dff/n5 ) );
  INV_X1 \product_reg/memory_57__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_57__dff/n7 ) );
  NAND2_X1 \product_reg/memory_57__dff/U3  ( .A1(\product_reg/n6 ), .A2(
        product_in[57]), .ZN(\product_reg/memory_57__dff/n6 ) );
  OAI21_X1 \product_reg/memory_57__dff/U2  ( .B1(\product_reg/n6 ), .B2(
        \product_reg/memory_57__dff/n5 ), .A(\product_reg/memory_57__dff/n6 ), 
        .ZN(\product_reg/memory_57__dff/n1 ) );
  DFFR_X1 \product_reg/memory_57__dff/q_reg  ( .D(
        \product_reg/memory_57__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_57__dff/n7 ), .Q(product_out[57]), .QN(
        \product_reg/memory_57__dff/n5 ) );
  INV_X1 \product_reg/memory_58__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_58__dff/n7 ) );
  NAND2_X1 \product_reg/memory_58__dff/U3  ( .A1(\product_reg/n6 ), .A2(
        product_in[58]), .ZN(\product_reg/memory_58__dff/n6 ) );
  OAI21_X1 \product_reg/memory_58__dff/U2  ( .B1(\product_reg/n6 ), .B2(
        \product_reg/memory_58__dff/n5 ), .A(\product_reg/memory_58__dff/n6 ), 
        .ZN(\product_reg/memory_58__dff/n1 ) );
  DFFR_X1 \product_reg/memory_58__dff/q_reg  ( .D(
        \product_reg/memory_58__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_58__dff/n7 ), .Q(product_out[58]), .QN(
        \product_reg/memory_58__dff/n5 ) );
  INV_X1 \product_reg/memory_59__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_59__dff/n7 ) );
  NAND2_X1 \product_reg/memory_59__dff/U3  ( .A1(\product_reg/n6 ), .A2(
        product_in[59]), .ZN(\product_reg/memory_59__dff/n6 ) );
  OAI21_X1 \product_reg/memory_59__dff/U2  ( .B1(\product_reg/n6 ), .B2(
        \product_reg/memory_59__dff/n5 ), .A(\product_reg/memory_59__dff/n6 ), 
        .ZN(\product_reg/memory_59__dff/n1 ) );
  DFFR_X1 \product_reg/memory_59__dff/q_reg  ( .D(
        \product_reg/memory_59__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_59__dff/n7 ), .Q(product_out[59]), .QN(
        \product_reg/memory_59__dff/n5 ) );
  INV_X1 \product_reg/memory_60__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_60__dff/n7 ) );
  NAND2_X1 \product_reg/memory_60__dff/U3  ( .A1(\product_reg/n7 ), .A2(
        product_in[60]), .ZN(\product_reg/memory_60__dff/n6 ) );
  OAI21_X1 \product_reg/memory_60__dff/U2  ( .B1(\product_reg/n7 ), .B2(
        \product_reg/memory_60__dff/n5 ), .A(\product_reg/memory_60__dff/n6 ), 
        .ZN(\product_reg/memory_60__dff/n1 ) );
  DFFR_X1 \product_reg/memory_60__dff/q_reg  ( .D(
        \product_reg/memory_60__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_60__dff/n7 ), .Q(product_out[60]), .QN(
        \product_reg/memory_60__dff/n5 ) );
  INV_X1 \product_reg/memory_61__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_61__dff/n7 ) );
  NAND2_X1 \product_reg/memory_61__dff/U3  ( .A1(\product_reg/n7 ), .A2(
        product_in[61]), .ZN(\product_reg/memory_61__dff/n6 ) );
  OAI21_X1 \product_reg/memory_61__dff/U2  ( .B1(\product_reg/n7 ), .B2(
        \product_reg/memory_61__dff/n5 ), .A(\product_reg/memory_61__dff/n6 ), 
        .ZN(\product_reg/memory_61__dff/n1 ) );
  DFFR_X1 \product_reg/memory_61__dff/q_reg  ( .D(
        \product_reg/memory_61__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_61__dff/n7 ), .Q(product_out[61]), .QN(
        \product_reg/memory_61__dff/n5 ) );
  NAND2_X1 \product_reg/memory_62__dff/U4  ( .A1(\product_reg/n7 ), .A2(n628), 
        .ZN(\product_reg/memory_62__dff/n6 ) );
  INV_X1 \product_reg/memory_62__dff/U3  ( .A(1'b0), .ZN(
        \product_reg/memory_62__dff/n7 ) );
  OAI21_X1 \product_reg/memory_62__dff/U2  ( .B1(\product_reg/n7 ), .B2(
        \product_reg/memory_62__dff/n5 ), .A(\product_reg/memory_62__dff/n6 ), 
        .ZN(\product_reg/memory_62__dff/n1 ) );
  DFFR_X1 \product_reg/memory_62__dff/q_reg  ( .D(
        \product_reg/memory_62__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_62__dff/n7 ), .Q(product_out[62]), .QN(
        \product_reg/memory_62__dff/n5 ) );
  NAND2_X1 \product_reg/memory_63__dff/U5  ( .A1(n631), .A2(\product_reg/n7 ), 
        .ZN(\product_reg/memory_63__dff/n7 ) );
  INV_X1 \product_reg/memory_63__dff/U4  ( .A(1'b0), .ZN(
        \product_reg/memory_63__dff/n8 ) );
  NAND2_X1 \product_reg/memory_63__dff/U3  ( .A1(
        \product_reg/memory_63__dff/n7 ), .A2(\product_reg/memory_63__dff/n5 ), 
        .ZN(\product_reg/memory_63__dff/n1 ) );
  OR2_X1 \product_reg/memory_63__dff/U2  ( .A1(\product_reg/n7 ), .A2(
        \product_reg/memory_63__dff/n6 ), .ZN(\product_reg/memory_63__dff/n5 )
         );
  DFFR_X1 \product_reg/memory_63__dff/q_reg  ( .D(
        \product_reg/memory_63__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_63__dff/n8 ), .Q(product_out[63]), .QN(
        \product_reg/memory_63__dff/n6 ) );
  OAI21_X1 \product_reg/memory_64__dff/U4  ( .B1(\product_reg/n7 ), .B2(
        \product_reg/memory_64__dff/n5 ), .A(\product_reg/memory_64__dff/n6 ), 
        .ZN(\product_reg/memory_64__dff/n1 ) );
  INV_X1 \product_reg/memory_64__dff/U3  ( .A(1'b0), .ZN(
        \product_reg/memory_64__dff/n7 ) );
  NAND2_X1 \product_reg/memory_64__dff/U2  ( .A1(\product_reg/n7 ), .A2(
        product_in[64]), .ZN(\product_reg/memory_64__dff/n6 ) );
  DFFR_X1 \product_reg/memory_64__dff/q_reg  ( .D(
        \product_reg/memory_64__dff/n1 ), .CK(clock), .RN(
        \product_reg/memory_64__dff/n7 ), .Q(product_out[64]), .QN(
        \product_reg/memory_64__dff/n5 ) );
endmodule

