
module multdiv ( data_operandA, data_operandB, ctrl_MULT, ctrl_DIV, clock, 
        data_result, data_exception, data_resultRDY, test_si1, test_so1, 
        test_si2, test_so2, test_si3, test_so3, test_se );
  input [31:0] data_operandA;
  input [31:0] data_operandB;
  output [31:0] data_result;
  input ctrl_MULT, ctrl_DIV, clock, test_si1, test_si2, test_si3, test_se;
  output data_exception, data_resultRDY, test_so1, test_so2, test_so3;
  wire   n187, n196, n197, n198, n209, n210, n212, n213, n214, n397, n625,
         \ctrl/op_div_int , \ctrl/mult_ready , \ctrl/op_mult_int ,
         \ctrl/counter/w7 , \ctrl/counter/w5 , \ctrl/cur_mult/n1 ,
         \ctrl/cur_div/n1 , \product_reg/memory_0__dff/n5 ,
         \product_reg/memory_1__dff/n8 , \product_reg/memory_1__dff/n1 ,
         \product_reg/memory_2__dff/n7 , \product_reg/memory_3__dff/n5 ,
         \product_reg/memory_3__dff/n1 , \product_reg/memory_4__dff/n5 ,
         \product_reg/memory_4__dff/n1 , \product_reg/memory_5__dff/n5 ,
         \product_reg/memory_5__dff/n1 , \product_reg/memory_6__dff/n5 ,
         \product_reg/memory_6__dff/n1 , \product_reg/memory_7__dff/n5 ,
         \product_reg/memory_7__dff/n1 , \product_reg/memory_8__dff/n5 ,
         \product_reg/memory_8__dff/n1 , \product_reg/memory_9__dff/n5 ,
         \product_reg/memory_9__dff/n1 , \product_reg/memory_10__dff/n5 ,
         \product_reg/memory_10__dff/n1 , \product_reg/memory_11__dff/n5 ,
         \product_reg/memory_11__dff/n1 , \product_reg/memory_12__dff/n5 ,
         \product_reg/memory_12__dff/n1 , \product_reg/memory_13__dff/n5 ,
         \product_reg/memory_13__dff/n1 , \product_reg/memory_14__dff/n5 ,
         \product_reg/memory_14__dff/n1 , \product_reg/memory_15__dff/n5 ,
         \product_reg/memory_15__dff/n1 , \product_reg/memory_16__dff/n5 ,
         \product_reg/memory_16__dff/n1 , \product_reg/memory_17__dff/n5 ,
         \product_reg/memory_17__dff/n1 , \product_reg/memory_18__dff/n5 ,
         \product_reg/memory_18__dff/n1 , \product_reg/memory_19__dff/n5 ,
         \product_reg/memory_19__dff/n1 , \product_reg/memory_20__dff/n5 ,
         \product_reg/memory_20__dff/n1 , \product_reg/memory_21__dff/n5 ,
         \product_reg/memory_21__dff/n1 , \product_reg/memory_22__dff/n5 ,
         \product_reg/memory_22__dff/n1 , \product_reg/memory_23__dff/n5 ,
         \product_reg/memory_23__dff/n1 , \product_reg/memory_24__dff/n5 ,
         \product_reg/memory_24__dff/n1 , \product_reg/memory_25__dff/n5 ,
         \product_reg/memory_25__dff/n1 , \product_reg/memory_26__dff/n5 ,
         \product_reg/memory_26__dff/n1 , \product_reg/memory_27__dff/n5 ,
         \product_reg/memory_27__dff/n1 , \product_reg/memory_28__dff/n5 ,
         \product_reg/memory_28__dff/n1 , \product_reg/memory_29__dff/n5 ,
         \product_reg/memory_29__dff/n1 , \product_reg/memory_30__dff/n5 ,
         \product_reg/memory_30__dff/n1 , \product_reg/memory_31__dff/n5 ,
         \product_reg/memory_31__dff/n1 , \product_reg/memory_32__dff/n1 ,
         \product_reg/memory_33__dff/n5 , \product_reg/memory_33__dff/n1 ,
         \product_reg/memory_34__dff/n5 , \product_reg/memory_34__dff/n1 ,
         \product_reg/memory_35__dff/n5 , \product_reg/memory_35__dff/n1 ,
         \product_reg/memory_36__dff/n5 , \product_reg/memory_36__dff/n1 ,
         \product_reg/memory_37__dff/n5 , \product_reg/memory_37__dff/n1 ,
         \product_reg/memory_38__dff/n5 , \product_reg/memory_38__dff/n1 ,
         \product_reg/memory_39__dff/n5 , \product_reg/memory_39__dff/n1 ,
         \product_reg/memory_40__dff/n5 , \product_reg/memory_40__dff/n1 ,
         \product_reg/memory_41__dff/n5 , \product_reg/memory_41__dff/n1 ,
         \product_reg/memory_42__dff/n5 , \product_reg/memory_42__dff/n1 ,
         \product_reg/memory_43__dff/n5 , \product_reg/memory_43__dff/n1 ,
         \product_reg/memory_44__dff/n5 , \product_reg/memory_44__dff/n1 ,
         \product_reg/memory_45__dff/n5 , \product_reg/memory_45__dff/n1 ,
         \product_reg/memory_46__dff/n5 , \product_reg/memory_46__dff/n1 ,
         \product_reg/memory_47__dff/n5 , \product_reg/memory_47__dff/n1 ,
         \product_reg/memory_48__dff/n5 , \product_reg/memory_48__dff/n1 ,
         \product_reg/memory_49__dff/n5 , \product_reg/memory_49__dff/n1 ,
         \product_reg/memory_50__dff/n5 , \product_reg/memory_50__dff/n1 ,
         \product_reg/memory_51__dff/n5 , \product_reg/memory_51__dff/n1 ,
         \product_reg/memory_52__dff/n5 , \product_reg/memory_52__dff/n1 ,
         \product_reg/memory_53__dff/n5 , \product_reg/memory_53__dff/n1 ,
         \product_reg/memory_54__dff/n5 , \product_reg/memory_54__dff/n1 ,
         \product_reg/memory_55__dff/n5 , \product_reg/memory_55__dff/n1 ,
         \product_reg/memory_56__dff/n5 , \product_reg/memory_56__dff/n1 ,
         \product_reg/memory_57__dff/n5 , \product_reg/memory_57__dff/n1 ,
         \product_reg/memory_58__dff/n5 , \product_reg/memory_58__dff/n1 ,
         \product_reg/memory_59__dff/n5 , \product_reg/memory_59__dff/n1 ,
         \product_reg/memory_60__dff/n5 , \product_reg/memory_60__dff/n1 ,
         \product_reg/memory_61__dff/n5 , \product_reg/memory_61__dff/n1 ,
         \product_reg/memory_62__dff/n5 , \product_reg/memory_62__dff/n1 ,
         \product_reg/memory_63__dff/n6 , \product_reg/memory_63__dff/n1 ,
         \product_reg/memory_64__dff/n5 , \product_reg/memory_64__dff/n1 , n65,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n112, n113, n115, n116, n117, n118, n119, n120, n122, n124,
         n126, n127, n128, n129, n130, n131, n132, n133, n135, n136, n137,
         n138, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n188, n189, n190, n191, n192, n193, n194,
         n195, n199, n200, n201, n202, n203, n204, n205, n206, n207, n211,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n473, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n704, n706, n708,
         n710, n713, n715, n717, n719, n721, n723, n725, n727, n729, n731,
         n733, n735, n737, n739, n741, n743, n745, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n758, n760, n761, n762, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1037, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071;
  wire   [64:0] product_out;
  wire   [31:0] adder_out;
  tri   [64:0] product_in;
  assign test_so2 = product_out[30];

  OAI22_X2 U1 ( .A1(data_resultRDY), .A2(n215), .B1(
        \product_reg/memory_9__dff/n5 ), .B2(n875), .ZN(
        \product_reg/memory_9__dff/n1 ) );
  INV_X4 U2 ( .A(product_in[9]), .ZN(n215) );
  OAI22_X2 U3 ( .A1(data_resultRDY), .A2(n217), .B1(
        \product_reg/memory_8__dff/n5 ), .B2(n873), .ZN(
        \product_reg/memory_8__dff/n1 ) );
  INV_X4 U4 ( .A(product_in[8]), .ZN(n217) );
  OAI22_X2 U5 ( .A1(data_resultRDY), .A2(n218), .B1(
        \product_reg/memory_7__dff/n5 ), .B2(n873), .ZN(
        \product_reg/memory_7__dff/n1 ) );
  INV_X4 U6 ( .A(product_in[7]), .ZN(n218) );
  OAI22_X2 U7 ( .A1(data_resultRDY), .A2(n219), .B1(
        \product_reg/memory_6__dff/n5 ), .B2(n873), .ZN(
        \product_reg/memory_6__dff/n1 ) );
  INV_X4 U8 ( .A(product_in[6]), .ZN(n219) );
  OAI22_X2 U9 ( .A1(data_resultRDY), .A2(n220), .B1(
        \product_reg/memory_64__dff/n5 ), .B2(n873), .ZN(
        \product_reg/memory_64__dff/n1 ) );
  INV_X4 U10 ( .A(product_in[64]), .ZN(n220) );
  OAI22_X2 U11 ( .A1(data_resultRDY), .A2(n221), .B1(
        \product_reg/memory_63__dff/n6 ), .B2(n873), .ZN(
        \product_reg/memory_63__dff/n1 ) );
  INV_X4 U12 ( .A(product_in[63]), .ZN(n221) );
  OAI22_X2 U13 ( .A1(data_resultRDY), .A2(n222), .B1(
        \product_reg/memory_62__dff/n5 ), .B2(n873), .ZN(
        \product_reg/memory_62__dff/n1 ) );
  OAI22_X2 U14 ( .A1(data_resultRDY), .A2(n223), .B1(
        \product_reg/memory_61__dff/n5 ), .B2(n873), .ZN(
        \product_reg/memory_61__dff/n1 ) );
  INV_X4 U15 ( .A(product_in[61]), .ZN(n223) );
  OAI22_X2 U16 ( .A1(data_resultRDY), .A2(n224), .B1(
        \product_reg/memory_60__dff/n5 ), .B2(n873), .ZN(
        \product_reg/memory_60__dff/n1 ) );
  INV_X4 U17 ( .A(product_in[60]), .ZN(n224) );
  OAI22_X2 U18 ( .A1(data_resultRDY), .A2(n225), .B1(
        \product_reg/memory_5__dff/n5 ), .B2(n873), .ZN(
        \product_reg/memory_5__dff/n1 ) );
  INV_X4 U19 ( .A(product_in[5]), .ZN(n225) );
  OAI22_X2 U20 ( .A1(n880), .A2(n226), .B1(\product_reg/memory_59__dff/n5 ), 
        .B2(n873), .ZN(\product_reg/memory_59__dff/n1 ) );
  INV_X4 U21 ( .A(product_in[59]), .ZN(n226) );
  OAI22_X2 U22 ( .A1(n880), .A2(n227), .B1(\product_reg/memory_58__dff/n5 ), 
        .B2(n873), .ZN(\product_reg/memory_58__dff/n1 ) );
  INV_X4 U23 ( .A(product_in[58]), .ZN(n227) );
  OAI22_X2 U24 ( .A1(n880), .A2(n228), .B1(\product_reg/memory_57__dff/n5 ), 
        .B2(n874), .ZN(\product_reg/memory_57__dff/n1 ) );
  INV_X4 U25 ( .A(product_in[57]), .ZN(n228) );
  OAI22_X2 U26 ( .A1(data_resultRDY), .A2(n229), .B1(
        \product_reg/memory_56__dff/n5 ), .B2(n874), .ZN(
        \product_reg/memory_56__dff/n1 ) );
  INV_X4 U27 ( .A(product_in[56]), .ZN(n229) );
  OAI22_X2 U28 ( .A1(data_resultRDY), .A2(n230), .B1(
        \product_reg/memory_55__dff/n5 ), .B2(n874), .ZN(
        \product_reg/memory_55__dff/n1 ) );
  INV_X4 U29 ( .A(product_in[55]), .ZN(n230) );
  OAI22_X2 U30 ( .A1(n880), .A2(n231), .B1(\product_reg/memory_54__dff/n5 ), 
        .B2(n874), .ZN(\product_reg/memory_54__dff/n1 ) );
  INV_X4 U31 ( .A(product_in[54]), .ZN(n231) );
  OAI22_X2 U32 ( .A1(data_resultRDY), .A2(n232), .B1(
        \product_reg/memory_53__dff/n5 ), .B2(n874), .ZN(
        \product_reg/memory_53__dff/n1 ) );
  INV_X4 U33 ( .A(product_in[53]), .ZN(n232) );
  OAI22_X2 U34 ( .A1(data_resultRDY), .A2(n233), .B1(
        \product_reg/memory_52__dff/n5 ), .B2(n874), .ZN(
        \product_reg/memory_52__dff/n1 ) );
  INV_X4 U35 ( .A(product_in[52]), .ZN(n233) );
  OAI22_X2 U36 ( .A1(data_resultRDY), .A2(n234), .B1(
        \product_reg/memory_51__dff/n5 ), .B2(n874), .ZN(
        \product_reg/memory_51__dff/n1 ) );
  INV_X4 U37 ( .A(product_in[51]), .ZN(n234) );
  OAI22_X2 U38 ( .A1(data_resultRDY), .A2(n235), .B1(
        \product_reg/memory_50__dff/n5 ), .B2(n874), .ZN(
        \product_reg/memory_50__dff/n1 ) );
  INV_X4 U39 ( .A(product_in[50]), .ZN(n235) );
  OAI22_X2 U40 ( .A1(data_resultRDY), .A2(n236), .B1(
        \product_reg/memory_4__dff/n5 ), .B2(n874), .ZN(
        \product_reg/memory_4__dff/n1 ) );
  INV_X4 U41 ( .A(product_in[4]), .ZN(n236) );
  OAI22_X2 U42 ( .A1(data_resultRDY), .A2(n237), .B1(
        \product_reg/memory_49__dff/n5 ), .B2(n874), .ZN(
        \product_reg/memory_49__dff/n1 ) );
  INV_X4 U43 ( .A(product_in[49]), .ZN(n237) );
  OAI22_X2 U44 ( .A1(n880), .A2(n238), .B1(\product_reg/memory_48__dff/n5 ), 
        .B2(n874), .ZN(\product_reg/memory_48__dff/n1 ) );
  INV_X4 U45 ( .A(product_in[48]), .ZN(n238) );
  OAI22_X2 U46 ( .A1(n880), .A2(n239), .B1(\product_reg/memory_47__dff/n5 ), 
        .B2(n874), .ZN(\product_reg/memory_47__dff/n1 ) );
  INV_X4 U47 ( .A(product_in[47]), .ZN(n239) );
  OAI22_X2 U48 ( .A1(n880), .A2(n240), .B1(\product_reg/memory_46__dff/n5 ), 
        .B2(n875), .ZN(\product_reg/memory_46__dff/n1 ) );
  INV_X4 U49 ( .A(product_in[46]), .ZN(n240) );
  OAI22_X2 U50 ( .A1(n880), .A2(n241), .B1(\product_reg/memory_45__dff/n5 ), 
        .B2(n875), .ZN(\product_reg/memory_45__dff/n1 ) );
  INV_X4 U51 ( .A(product_in[45]), .ZN(n241) );
  OAI22_X2 U52 ( .A1(n880), .A2(n242), .B1(\product_reg/memory_44__dff/n5 ), 
        .B2(n875), .ZN(\product_reg/memory_44__dff/n1 ) );
  INV_X4 U53 ( .A(product_in[44]), .ZN(n242) );
  OAI22_X2 U54 ( .A1(n880), .A2(n243), .B1(\product_reg/memory_43__dff/n5 ), 
        .B2(n875), .ZN(\product_reg/memory_43__dff/n1 ) );
  INV_X4 U55 ( .A(product_in[43]), .ZN(n243) );
  OAI22_X2 U56 ( .A1(n880), .A2(n244), .B1(\product_reg/memory_42__dff/n5 ), 
        .B2(n875), .ZN(\product_reg/memory_42__dff/n1 ) );
  INV_X4 U57 ( .A(product_in[42]), .ZN(n244) );
  OAI22_X2 U58 ( .A1(n880), .A2(n245), .B1(\product_reg/memory_41__dff/n5 ), 
        .B2(n875), .ZN(\product_reg/memory_41__dff/n1 ) );
  INV_X4 U59 ( .A(product_in[41]), .ZN(n245) );
  OAI22_X2 U60 ( .A1(n880), .A2(n246), .B1(\product_reg/memory_40__dff/n5 ), 
        .B2(n875), .ZN(\product_reg/memory_40__dff/n1 ) );
  INV_X4 U61 ( .A(product_in[40]), .ZN(n246) );
  OAI22_X2 U62 ( .A1(n880), .A2(n247), .B1(\product_reg/memory_3__dff/n5 ), 
        .B2(n875), .ZN(\product_reg/memory_3__dff/n1 ) );
  INV_X4 U63 ( .A(product_in[3]), .ZN(n247) );
  OAI22_X2 U64 ( .A1(n879), .A2(n248), .B1(\product_reg/memory_39__dff/n5 ), 
        .B2(n875), .ZN(\product_reg/memory_39__dff/n1 ) );
  INV_X4 U65 ( .A(product_in[39]), .ZN(n248) );
  OAI22_X2 U66 ( .A1(n879), .A2(n249), .B1(\product_reg/memory_38__dff/n5 ), 
        .B2(n875), .ZN(\product_reg/memory_38__dff/n1 ) );
  INV_X4 U67 ( .A(product_in[38]), .ZN(n249) );
  OAI22_X2 U68 ( .A1(n879), .A2(n250), .B1(\product_reg/memory_37__dff/n5 ), 
        .B2(n875), .ZN(\product_reg/memory_37__dff/n1 ) );
  INV_X4 U69 ( .A(product_in[37]), .ZN(n250) );
  OAI22_X2 U70 ( .A1(n879), .A2(n251), .B1(\product_reg/memory_36__dff/n5 ), 
        .B2(n876), .ZN(\product_reg/memory_36__dff/n1 ) );
  INV_X4 U71 ( .A(product_in[36]), .ZN(n251) );
  OAI22_X2 U72 ( .A1(n880), .A2(n252), .B1(\product_reg/memory_35__dff/n5 ), 
        .B2(n876), .ZN(\product_reg/memory_35__dff/n1 ) );
  INV_X4 U73 ( .A(product_in[35]), .ZN(n252) );
  OAI22_X2 U74 ( .A1(n880), .A2(n253), .B1(\product_reg/memory_34__dff/n5 ), 
        .B2(n876), .ZN(\product_reg/memory_34__dff/n1 ) );
  INV_X4 U75 ( .A(product_in[34]), .ZN(n253) );
  OAI22_X2 U76 ( .A1(n880), .A2(n254), .B1(\product_reg/memory_33__dff/n5 ), 
        .B2(n876), .ZN(\product_reg/memory_33__dff/n1 ) );
  INV_X4 U77 ( .A(product_in[33]), .ZN(n254) );
  OAI22_X2 U78 ( .A1(n880), .A2(n255), .B1(n878), .B2(n135), .ZN(
        \product_reg/memory_32__dff/n1 ) );
  INV_X4 U79 ( .A(product_in[32]), .ZN(n255) );
  OAI22_X2 U80 ( .A1(n880), .A2(n256), .B1(\product_reg/memory_31__dff/n5 ), 
        .B2(n876), .ZN(\product_reg/memory_31__dff/n1 ) );
  INV_X4 U81 ( .A(product_in[31]), .ZN(n256) );
  OAI22_X2 U82 ( .A1(n880), .A2(n257), .B1(\product_reg/memory_30__dff/n5 ), 
        .B2(n876), .ZN(\product_reg/memory_30__dff/n1 ) );
  INV_X4 U83 ( .A(product_in[30]), .ZN(n257) );
  OAI22_X2 U84 ( .A1(n880), .A2(n258), .B1(\product_reg/memory_29__dff/n5 ), 
        .B2(n876), .ZN(\product_reg/memory_29__dff/n1 ) );
  INV_X4 U85 ( .A(product_in[29]), .ZN(n258) );
  OAI22_X2 U86 ( .A1(n879), .A2(n259), .B1(\product_reg/memory_28__dff/n5 ), 
        .B2(n876), .ZN(\product_reg/memory_28__dff/n1 ) );
  INV_X4 U87 ( .A(product_in[28]), .ZN(n259) );
  OAI22_X2 U88 ( .A1(n879), .A2(n260), .B1(\product_reg/memory_27__dff/n5 ), 
        .B2(n876), .ZN(\product_reg/memory_27__dff/n1 ) );
  INV_X4 U89 ( .A(product_in[27]), .ZN(n260) );
  OAI22_X2 U90 ( .A1(n879), .A2(n261), .B1(\product_reg/memory_26__dff/n5 ), 
        .B2(n876), .ZN(\product_reg/memory_26__dff/n1 ) );
  INV_X4 U91 ( .A(product_in[26]), .ZN(n261) );
  OAI22_X2 U92 ( .A1(n879), .A2(n262), .B1(\product_reg/memory_25__dff/n5 ), 
        .B2(n876), .ZN(\product_reg/memory_25__dff/n1 ) );
  INV_X4 U93 ( .A(product_in[25]), .ZN(n262) );
  OAI22_X2 U94 ( .A1(n879), .A2(n263), .B1(\product_reg/memory_24__dff/n5 ), 
        .B2(n876), .ZN(\product_reg/memory_24__dff/n1 ) );
  INV_X4 U95 ( .A(product_in[24]), .ZN(n263) );
  OAI22_X2 U96 ( .A1(n879), .A2(n264), .B1(\product_reg/memory_23__dff/n5 ), 
        .B2(n877), .ZN(\product_reg/memory_23__dff/n1 ) );
  INV_X4 U97 ( .A(product_in[23]), .ZN(n264) );
  OAI22_X2 U98 ( .A1(n879), .A2(n265), .B1(\product_reg/memory_22__dff/n5 ), 
        .B2(n877), .ZN(\product_reg/memory_22__dff/n1 ) );
  INV_X4 U99 ( .A(product_in[22]), .ZN(n265) );
  OAI22_X2 U100 ( .A1(n879), .A2(n266), .B1(\product_reg/memory_21__dff/n5 ), 
        .B2(n877), .ZN(\product_reg/memory_21__dff/n1 ) );
  INV_X4 U101 ( .A(product_in[21]), .ZN(n266) );
  OAI22_X2 U102 ( .A1(n879), .A2(n267), .B1(\product_reg/memory_20__dff/n5 ), 
        .B2(n877), .ZN(\product_reg/memory_20__dff/n1 ) );
  INV_X4 U103 ( .A(product_in[20]), .ZN(n267) );
  OAI22_X2 U104 ( .A1(n879), .A2(n268), .B1(\product_reg/memory_1__dff/n8 ), 
        .B2(n877), .ZN(\product_reg/memory_1__dff/n1 ) );
  INV_X4 U105 ( .A(product_in[1]), .ZN(n268) );
  OAI22_X2 U106 ( .A1(n879), .A2(n269), .B1(\product_reg/memory_19__dff/n5 ), 
        .B2(n877), .ZN(\product_reg/memory_19__dff/n1 ) );
  INV_X4 U107 ( .A(product_in[19]), .ZN(n269) );
  OAI22_X2 U108 ( .A1(n879), .A2(n270), .B1(\product_reg/memory_18__dff/n5 ), 
        .B2(n877), .ZN(\product_reg/memory_18__dff/n1 ) );
  INV_X4 U109 ( .A(product_in[18]), .ZN(n270) );
  OAI22_X2 U110 ( .A1(n880), .A2(n271), .B1(\product_reg/memory_17__dff/n5 ), 
        .B2(n877), .ZN(\product_reg/memory_17__dff/n1 ) );
  INV_X4 U111 ( .A(product_in[17]), .ZN(n271) );
  OAI22_X2 U112 ( .A1(n879), .A2(n272), .B1(\product_reg/memory_16__dff/n5 ), 
        .B2(n877), .ZN(\product_reg/memory_16__dff/n1 ) );
  INV_X4 U113 ( .A(product_in[16]), .ZN(n272) );
  OAI22_X2 U114 ( .A1(n879), .A2(n273), .B1(\product_reg/memory_15__dff/n5 ), 
        .B2(n877), .ZN(\product_reg/memory_15__dff/n1 ) );
  INV_X4 U115 ( .A(product_in[15]), .ZN(n273) );
  OAI22_X2 U116 ( .A1(n879), .A2(n274), .B1(\product_reg/memory_14__dff/n5 ), 
        .B2(n877), .ZN(\product_reg/memory_14__dff/n1 ) );
  INV_X4 U117 ( .A(product_in[14]), .ZN(n274) );
  OAI22_X2 U118 ( .A1(n879), .A2(n275), .B1(\product_reg/memory_13__dff/n5 ), 
        .B2(n877), .ZN(\product_reg/memory_13__dff/n1 ) );
  INV_X4 U119 ( .A(product_in[13]), .ZN(n275) );
  OAI22_X2 U120 ( .A1(n879), .A2(n276), .B1(\product_reg/memory_12__dff/n5 ), 
        .B2(n878), .ZN(\product_reg/memory_12__dff/n1 ) );
  INV_X4 U121 ( .A(product_in[12]), .ZN(n276) );
  OAI22_X2 U122 ( .A1(n879), .A2(n277), .B1(\product_reg/memory_11__dff/n5 ), 
        .B2(n878), .ZN(\product_reg/memory_11__dff/n1 ) );
  INV_X4 U123 ( .A(product_in[11]), .ZN(n277) );
  OAI22_X2 U124 ( .A1(n879), .A2(n278), .B1(\product_reg/memory_10__dff/n5 ), 
        .B2(n878), .ZN(\product_reg/memory_10__dff/n1 ) );
  INV_X4 U125 ( .A(product_in[10]), .ZN(n278) );
  AOI22_X2 U126 ( .A1(n873), .A2(product_in[0]), .B1(n118), .B2(data_resultRDY), .ZN(n279) );
  OAI22_X2 U128 ( .A1(\product_reg/memory_30__dff/n5 ), .A2(n869), .B1(n280), 
        .B2(n871), .ZN(data_result[29]) );
  OAI22_X2 U129 ( .A1(data_operandA[31]), .A2(n141), .B1(n898), .B2(n280), 
        .ZN(n704) );
  XNOR2_X2 U130 ( .A(n282), .B(n283), .ZN(n280) );
  OR2_X2 U131 ( .A1(n284), .A2(n285), .ZN(n282) );
  OAI22_X2 U132 ( .A1(\product_reg/memory_29__dff/n5 ), .A2(n869), .B1(n871), 
        .B2(n286), .ZN(data_result[28]) );
  OAI22_X2 U133 ( .A1(data_operandA[31]), .A2(n142), .B1(n897), .B2(n286), 
        .ZN(n706) );
  XNOR2_X2 U134 ( .A(n284), .B(n285), .ZN(n286) );
  OAI22_X2 U135 ( .A1(\product_reg/memory_25__dff/n5 ), .A2(n869), .B1(n287), 
        .B2(n871), .ZN(data_result[24]) );
  OAI22_X2 U136 ( .A1(data_operandA[31]), .A2(n146), .B1(n287), .B2(n897), 
        .ZN(n708) );
  XNOR2_X2 U137 ( .A(n288), .B(n289), .ZN(n287) );
  OAI22_X2 U138 ( .A1(\product_reg/memory_27__dff/n5 ), .A2(n869), .B1(n871), 
        .B2(n290), .ZN(data_result[26]) );
  OAI22_X2 U139 ( .A1(data_operandA[31]), .A2(n144), .B1(n897), .B2(n290), 
        .ZN(n710) );
  XNOR2_X2 U140 ( .A(n291), .B(n292), .ZN(n290) );
  OAI22_X2 U141 ( .A1(\product_reg/memory_31__dff/n5 ), .A2(n869), .B1(n871), 
        .B2(n293), .ZN(data_result[30]) );
  OAI22_X2 U142 ( .A1(\product_reg/memory_28__dff/n5 ), .A2(n869), .B1(n871), 
        .B2(n294), .ZN(data_result[27]) );
  OAI22_X2 U143 ( .A1(data_operandA[31]), .A2(n143), .B1(n897), .B2(n294), 
        .ZN(n713) );
  XNOR2_X2 U144 ( .A(n295), .B(n296), .ZN(n294) );
  OR2_X2 U145 ( .A1(n291), .A2(n292), .ZN(n295) );
  OAI22_X2 U146 ( .A1(\product_reg/memory_26__dff/n5 ), .A2(n869), .B1(n871), 
        .B2(n297), .ZN(data_result[25]) );
  OAI22_X2 U147 ( .A1(data_operandA[31]), .A2(n145), .B1(n897), .B2(n297), 
        .ZN(n715) );
  XNOR2_X2 U148 ( .A(n298), .B(n299), .ZN(n297) );
  OR2_X2 U149 ( .A1(n289), .A2(n288), .ZN(n298) );
  OAI22_X2 U150 ( .A1(\product_reg/memory_24__dff/n5 ), .A2(n869), .B1(n871), 
        .B2(n300), .ZN(data_result[23]) );
  OAI22_X2 U151 ( .A1(data_operandA[31]), .A2(n147), .B1(n897), .B2(n300), 
        .ZN(n717) );
  XNOR2_X2 U152 ( .A(n301), .B(n302), .ZN(n300) );
  NAND2_X2 U153 ( .A1(n303), .A2(n133), .ZN(n301) );
  OAI22_X2 U154 ( .A1(data_operandA[31]), .A2(n151), .B1(n897), .B2(n305), 
        .ZN(n719) );
  OAI22_X2 U155 ( .A1(data_operandA[31]), .A2(n152), .B1(n897), .B2(n306), 
        .ZN(n721) );
  OAI22_X2 U156 ( .A1(data_operandA[31]), .A2(n153), .B1(n897), .B2(n307), 
        .ZN(n723) );
  OAI22_X2 U157 ( .A1(data_operandA[31]), .A2(n154), .B1(n897), .B2(n308), 
        .ZN(n725) );
  OAI22_X2 U158 ( .A1(data_operandA[31]), .A2(n155), .B1(n897), .B2(n309), 
        .ZN(n727) );
  OAI22_X2 U159 ( .A1(data_operandA[31]), .A2(n156), .B1(n897), .B2(n310), 
        .ZN(n729) );
  OAI22_X2 U160 ( .A1(data_operandA[31]), .A2(n157), .B1(n898), .B2(n311), 
        .ZN(n731) );
  OAI22_X2 U161 ( .A1(data_operandA[31]), .A2(n159), .B1(n898), .B2(n312), 
        .ZN(n733) );
  OAI22_X2 U162 ( .A1(data_operandA[31]), .A2(n160), .B1(n898), .B2(n313), 
        .ZN(n735) );
  OAI22_X2 U163 ( .A1(data_operandA[31]), .A2(n158), .B1(n898), .B2(n314), 
        .ZN(n737) );
  OAI22_X2 U164 ( .A1(\product_reg/memory_3__dff/n5 ), .A2(n869), .B1(n871), 
        .B2(n315), .ZN(data_result[2]) );
  OAI22_X2 U165 ( .A1(data_operandA[31]), .A2(n168), .B1(n898), .B2(n315), 
        .ZN(n739) );
  XNOR2_X2 U166 ( .A(n316), .B(n317), .ZN(n315) );
  OAI22_X2 U167 ( .A1(\product_reg/memory_5__dff/n5 ), .A2(n870), .B1(n871), 
        .B2(n318), .ZN(data_result[4]) );
  OAI22_X2 U168 ( .A1(data_operandA[31]), .A2(n166), .B1(n898), .B2(n318), 
        .ZN(n741) );
  XNOR2_X2 U169 ( .A(n319), .B(n320), .ZN(n318) );
  OAI22_X2 U170 ( .A1(\product_reg/memory_4__dff/n5 ), .A2(n870), .B1(n871), 
        .B2(n321), .ZN(data_result[3]) );
  OAI22_X2 U171 ( .A1(data_operandA[31]), .A2(n167), .B1(n898), .B2(n321), 
        .ZN(n743) );
  XOR2_X2 U172 ( .A(n322), .B(n323), .Z(n321) );
  OAI22_X2 U173 ( .A1(\product_reg/memory_2__dff/n7 ), .A2(n870), .B1(n324), 
        .B2(n871), .ZN(data_result[1]) );
  OAI22_X2 U174 ( .A1(data_operandA[31]), .A2(n169), .B1(n324), .B2(n897), 
        .ZN(n745) );
  XNOR2_X2 U175 ( .A(n325), .B(n326), .ZN(n324) );
  OAI22_X2 U176 ( .A1(data_operandA[31]), .A2(n170), .B1(n325), .B2(n897), 
        .ZN(n747) );
  OAI22_X2 U177 ( .A1(product_in[2]), .A2(data_resultRDY), .B1(n878), .B2(
        product_out[2]), .ZN(n755) );
  OAI22_X2 U178 ( .A1(data_operandA[31]), .A2(n140), .B1(n898), .B2(n293), 
        .ZN(n397) );
  XNOR2_X2 U179 ( .A(n327), .B(n328), .ZN(n293) );
  OAI22_X2 U180 ( .A1(data_operandA[31]), .A2(n165), .B1(n898), .B2(n329), 
        .ZN(n214) );
  OAI22_X2 U181 ( .A1(data_operandA[31]), .A2(n164), .B1(n898), .B2(n330), 
        .ZN(n213) );
  OAI22_X2 U182 ( .A1(data_operandA[31]), .A2(n163), .B1(n898), .B2(n331), 
        .ZN(n212) );
  OAI22_X2 U183 ( .A1(data_operandA[31]), .A2(n162), .B1(n898), .B2(n332), 
        .ZN(n210) );
  OAI22_X2 U184 ( .A1(data_operandA[31]), .A2(n161), .B1(n898), .B2(n333), 
        .ZN(n209) );
  OAI22_X2 U185 ( .A1(data_operandA[31]), .A2(n150), .B1(n898), .B2(n334), 
        .ZN(n198) );
  OAI22_X2 U186 ( .A1(data_operandA[31]), .A2(n149), .B1(n898), .B2(n335), 
        .ZN(n197) );
  OAI22_X2 U187 ( .A1(data_operandA[31]), .A2(n148), .B1(n897), .B2(n336), 
        .ZN(n196) );
  INV_X4 U190 ( .A(product_in[62]), .ZN(n222) );
  OAI22_X2 U191 ( .A1(\product_reg/memory_10__dff/n5 ), .A2(n870), .B1(n871), 
        .B2(n333), .ZN(data_result[9]) );
  XNOR2_X2 U192 ( .A(n338), .B(n339), .ZN(n333) );
  OAI22_X2 U193 ( .A1(\product_reg/memory_9__dff/n5 ), .A2(n870), .B1(n871), 
        .B2(n332), .ZN(data_result[8]) );
  XNOR2_X2 U194 ( .A(n340), .B(n341), .ZN(n332) );
  OAI22_X2 U195 ( .A1(\product_reg/memory_8__dff/n5 ), .A2(n870), .B1(n871), 
        .B2(n331), .ZN(data_result[7]) );
  XNOR2_X2 U196 ( .A(n342), .B(n343), .ZN(n331) );
  OAI22_X2 U197 ( .A1(\product_reg/memory_7__dff/n5 ), .A2(n870), .B1(n871), 
        .B2(n330), .ZN(data_result[6]) );
  XOR2_X2 U198 ( .A(n344), .B(n124), .Z(n330) );
  NAND2_X2 U199 ( .A1(n345), .A2(n346), .ZN(n344) );
  OAI22_X2 U200 ( .A1(\product_reg/memory_6__dff/n5 ), .A2(n870), .B1(n871), 
        .B2(n329), .ZN(data_result[5]) );
  XNOR2_X2 U201 ( .A(n346), .B(n345), .ZN(n329) );
  OAI22_X2 U202 ( .A1(\product_reg/memory_23__dff/n5 ), .A2(n870), .B1(n871), 
        .B2(n336), .ZN(data_result[22]) );
  XOR2_X2 U203 ( .A(n304), .B(n303), .Z(n336) );
  OAI22_X2 U205 ( .A1(\product_reg/memory_22__dff/n5 ), .A2(n870), .B1(n871), 
        .B2(n335), .ZN(data_result[21]) );
  XOR2_X2 U206 ( .A(n347), .B(n350), .Z(n335) );
  OAI22_X2 U208 ( .A1(\product_reg/memory_21__dff/n5 ), .A2(n870), .B1(n871), 
        .B2(n334), .ZN(data_result[20]) );
  XNOR2_X2 U209 ( .A(n349), .B(n348), .ZN(n334) );
  OAI22_X2 U211 ( .A1(n352), .A2(n762), .B1(n702), .B2(n353), .ZN(
        data_exception) );
  NOR4_X2 U213 ( .A1(n357), .A2(n358), .A3(n359), .A4(n360), .ZN(n355) );
  NAND4_X2 U214 ( .A1(n178), .A2(n177), .A3(n176), .A4(n175), .ZN(n360) );
  NAND4_X2 U215 ( .A1(n174), .A2(n173), .A3(n204), .A4(n172), .ZN(n359) );
  NAND4_X2 U216 ( .A1(n171), .A2(n203), .A3(n202), .A4(n201), .ZN(n358) );
  NAND4_X2 U217 ( .A1(n200), .A2(n199), .A3(n195), .A4(n194), .ZN(n357) );
  NOR4_X2 U218 ( .A1(n361), .A2(n362), .A3(n363), .A4(n364), .ZN(n354) );
  NAND4_X2 U219 ( .A1(n206), .A2(n193), .A3(n192), .A4(n191), .ZN(n364) );
  NAND4_X2 U220 ( .A1(n190), .A2(n189), .A3(n188), .A4(n186), .ZN(n363) );
  NAND4_X2 U221 ( .A1(n185), .A2(n184), .A3(n183), .A4(n205), .ZN(n362) );
  NAND4_X2 U222 ( .A1(n182), .A2(n181), .A3(n180), .A4(n179), .ZN(n361) );
  NAND4_X2 U224 ( .A1(n369), .A2(n370), .A3(n371), .A4(n372), .ZN(n368) );
  NOR4_X2 U225 ( .A1(n373), .A2(n374), .A3(n375), .A4(n376), .ZN(n372) );
  OR4_X2 U226 ( .A1(n135), .A2(\product_reg/memory_33__dff/n5 ), .A3(
        \product_reg/memory_34__dff/n5 ), .A4(\product_reg/memory_35__dff/n5 ), 
        .ZN(n376) );
  OR4_X2 U227 ( .A1(\product_reg/memory_36__dff/n5 ), .A2(
        \product_reg/memory_37__dff/n5 ), .A3(\product_reg/memory_38__dff/n5 ), 
        .A4(\product_reg/memory_39__dff/n5 ), .ZN(n375) );
  OR4_X2 U228 ( .A1(\product_reg/memory_40__dff/n5 ), .A2(
        \product_reg/memory_41__dff/n5 ), .A3(\product_reg/memory_42__dff/n5 ), 
        .A4(\product_reg/memory_43__dff/n5 ), .ZN(n374) );
  OR4_X2 U229 ( .A1(\product_reg/memory_44__dff/n5 ), .A2(
        \product_reg/memory_45__dff/n5 ), .A3(\product_reg/memory_46__dff/n5 ), 
        .A4(\product_reg/memory_47__dff/n5 ), .ZN(n373) );
  NOR4_X2 U230 ( .A1(n377), .A2(n378), .A3(\product_reg/memory_61__dff/n5 ), 
        .A4(\product_reg/memory_60__dff/n5 ), .ZN(n371) );
  OR3_X2 U231 ( .A1(\product_reg/memory_63__dff/n6 ), .A2(
        \product_reg/memory_64__dff/n5 ), .A3(\product_reg/memory_62__dff/n5 ), 
        .ZN(n378) );
  OR4_X2 U232 ( .A1(\product_reg/memory_56__dff/n5 ), .A2(
        \product_reg/memory_57__dff/n5 ), .A3(\product_reg/memory_58__dff/n5 ), 
        .A4(\product_reg/memory_59__dff/n5 ), .ZN(n377) );
  NOR4_X2 U233 ( .A1(\product_reg/memory_55__dff/n5 ), .A2(
        \product_reg/memory_54__dff/n5 ), .A3(\product_reg/memory_53__dff/n5 ), 
        .A4(\product_reg/memory_52__dff/n5 ), .ZN(n370) );
  NOR4_X2 U234 ( .A1(\product_reg/memory_51__dff/n5 ), .A2(
        \product_reg/memory_50__dff/n5 ), .A3(\product_reg/memory_49__dff/n5 ), 
        .A4(\product_reg/memory_48__dff/n5 ), .ZN(n369) );
  NAND4_X2 U235 ( .A1(n379), .A2(n380), .A3(n381), .A4(n382), .ZN(n367) );
  NOR4_X2 U236 ( .A1(n383), .A2(n384), .A3(n385), .A4(n386), .ZN(n382) );
  NAND4_X2 U237 ( .A1(\product_reg/memory_64__dff/n5 ), .A2(
        \product_reg/memory_61__dff/n5 ), .A3(\product_reg/memory_56__dff/n5 ), 
        .A4(\product_reg/memory_53__dff/n5 ), .ZN(n386) );
  NAND4_X2 U238 ( .A1(\product_reg/memory_48__dff/n5 ), .A2(
        \product_reg/memory_45__dff/n5 ), .A3(\product_reg/memory_40__dff/n5 ), 
        .A4(\product_reg/memory_37__dff/n5 ), .ZN(n385) );
  NAND4_X2 U239 ( .A1(\product_reg/memory_36__dff/n5 ), .A2(
        \product_reg/memory_35__dff/n5 ), .A3(\product_reg/memory_34__dff/n5 ), 
        .A4(\product_reg/memory_33__dff/n5 ), .ZN(n384) );
  NAND4_X2 U240 ( .A1(\product_reg/memory_60__dff/n5 ), .A2(
        \product_reg/memory_59__dff/n5 ), .A3(\product_reg/memory_58__dff/n5 ), 
        .A4(\product_reg/memory_57__dff/n5 ), .ZN(n383) );
  NOR4_X2 U241 ( .A1(n387), .A2(n388), .A3(n136), .A4(n137), .ZN(n381) );
  NAND4_X2 U243 ( .A1(\product_reg/memory_47__dff/n5 ), .A2(
        \product_reg/memory_46__dff/n5 ), .A3(\product_reg/memory_50__dff/n5 ), 
        .A4(\product_reg/memory_49__dff/n5 ), .ZN(n387) );
  AND4_X2 U244 ( .A1(\product_reg/memory_41__dff/n5 ), .A2(
        \product_reg/memory_42__dff/n5 ), .A3(\product_reg/memory_38__dff/n5 ), 
        .A4(\product_reg/memory_39__dff/n5 ), .ZN(n380) );
  AND4_X2 U245 ( .A1(\product_reg/memory_43__dff/n5 ), .A2(
        \product_reg/memory_44__dff/n5 ), .A3(\product_reg/memory_51__dff/n5 ), 
        .A4(\product_reg/memory_52__dff/n5 ), .ZN(n379) );
  NOR4_X2 U247 ( .A1(n390), .A2(n391), .A3(n392), .A4(n393), .ZN(n389) );
  NAND4_X2 U248 ( .A1(\product_reg/memory_22__dff/n5 ), .A2(
        \product_reg/memory_21__dff/n5 ), .A3(\product_reg/memory_23__dff/n5 ), 
        .A4(\product_reg/memory_24__dff/n5 ), .ZN(n393) );
  NAND4_X2 U249 ( .A1(\product_reg/memory_8__dff/n5 ), .A2(
        \product_reg/memory_7__dff/n5 ), .A3(\product_reg/memory_4__dff/n5 ), 
        .A4(\product_reg/memory_3__dff/n5 ), .ZN(n392) );
  NAND4_X2 U250 ( .A1(\product_reg/memory_31__dff/n5 ), .A2(
        \product_reg/memory_29__dff/n5 ), .A3(\product_reg/memory_2__dff/n7 ), 
        .A4(n394), .ZN(n391) );
  AND4_X2 U251 ( .A1(\product_reg/memory_25__dff/n5 ), .A2(
        \product_reg/memory_26__dff/n5 ), .A3(\product_reg/memory_27__dff/n5 ), 
        .A4(\product_reg/memory_28__dff/n5 ), .ZN(n394) );
  NAND4_X2 U252 ( .A1(n395), .A2(n396), .A3(n398), .A4(n399), .ZN(n390) );
  NOR4_X2 U253 ( .A1(data_result[19]), .A2(data_result[18]), .A3(
        data_result[17]), .A4(data_result[16]), .ZN(n399) );
  OAI22_X2 U254 ( .A1(\product_reg/memory_17__dff/n5 ), .A2(n870), .B1(n872), 
        .B2(n308), .ZN(data_result[16]) );
  XNOR2_X2 U255 ( .A(n400), .B(n401), .ZN(n308) );
  OAI22_X2 U256 ( .A1(\product_reg/memory_18__dff/n5 ), .A2(n869), .B1(n872), 
        .B2(n307), .ZN(data_result[17]) );
  XOR2_X2 U257 ( .A(n402), .B(n403), .Z(n307) );
  OAI22_X2 U259 ( .A1(\product_reg/memory_19__dff/n5 ), .A2(n834), .B1(n872), 
        .B2(n306), .ZN(data_result[18]) );
  XOR2_X2 U260 ( .A(n404), .B(n351), .Z(n306) );
  OAI22_X2 U261 ( .A1(\product_reg/memory_20__dff/n5 ), .A2(n834), .B1(n872), 
        .B2(n305), .ZN(data_result[19]) );
  XOR2_X2 U262 ( .A(n405), .B(n131), .Z(n305) );
  NAND2_X2 U263 ( .A1(n351), .A2(n130), .ZN(n405) );
  NOR4_X2 U265 ( .A1(data_result[15]), .A2(data_result[14]), .A3(
        data_result[13]), .A4(data_result[11]), .ZN(n398) );
  OAI22_X2 U266 ( .A1(\product_reg/memory_12__dff/n5 ), .A2(n834), .B1(n872), 
        .B2(n312), .ZN(data_result[11]) );
  XOR2_X2 U267 ( .A(n406), .B(n127), .Z(n312) );
  NAND2_X2 U268 ( .A1(n407), .A2(n126), .ZN(n406) );
  OAI22_X2 U269 ( .A1(\product_reg/memory_14__dff/n5 ), .A2(n834), .B1(n872), 
        .B2(n311), .ZN(data_result[13]) );
  XOR2_X2 U270 ( .A(n408), .B(n409), .Z(n311) );
  OAI22_X2 U272 ( .A1(\product_reg/memory_15__dff/n5 ), .A2(n834), .B1(n872), 
        .B2(n310), .ZN(data_result[14]) );
  XOR2_X2 U273 ( .A(n412), .B(n413), .Z(n310) );
  OAI22_X2 U274 ( .A1(\product_reg/memory_16__dff/n5 ), .A2(n834), .B1(n872), 
        .B2(n309), .ZN(data_result[15]) );
  XOR2_X2 U275 ( .A(n414), .B(n129), .Z(n309) );
  NAND2_X2 U276 ( .A1(n413), .A2(n128), .ZN(n414) );
  NOR4_X2 U277 ( .A1(data_result[10]), .A2(data_result[12]), .A3(
        data_result[0]), .A4(product_out[30]), .ZN(n396) );
  OAI22_X2 U278 ( .A1(\product_reg/memory_1__dff/n8 ), .A2(n834), .B1(n325), 
        .B2(n871), .ZN(data_result[0]) );
  OAI22_X2 U279 ( .A1(\product_reg/memory_13__dff/n5 ), .A2(n834), .B1(n872), 
        .B2(n314), .ZN(data_result[12]) );
  XNOR2_X2 U280 ( .A(n411), .B(n410), .ZN(n314) );
  OAI22_X2 U281 ( .A1(\product_reg/memory_11__dff/n5 ), .A2(n834), .B1(n871), 
        .B2(n313), .ZN(data_result[10]) );
  XOR2_X2 U282 ( .A(n415), .B(n407), .Z(n313) );
  AND4_X2 U283 ( .A1(\product_reg/memory_10__dff/n5 ), .A2(
        \product_reg/memory_9__dff/n5 ), .A3(\product_reg/memory_6__dff/n5 ), 
        .A4(\product_reg/memory_5__dff/n5 ), .ZN(n395) );
  OAI22_X2 U284 ( .A1(n869), .A2(n135), .B1(n337), .B2(n872), .ZN(
        data_result[31]) );
  OAI22_X2 U288 ( .A1(data_operandA[31]), .A2(n896), .B1(product_out[32]), 
        .B2(ctrl_DIV), .ZN(n417) );
  AOI22_X2 U289 ( .A1(n140), .A2(ctrl_DIV), .B1(n896), .B2(
        \product_reg/memory_31__dff/n5 ), .ZN(n328) );
  OR3_X2 U290 ( .A1(n285), .A2(n283), .A3(n284), .ZN(n327) );
  OR3_X2 U291 ( .A1(n296), .A2(n292), .A3(n291), .ZN(n284) );
  OR3_X2 U292 ( .A1(n289), .A2(n288), .A3(n299), .ZN(n291) );
  AOI22_X2 U293 ( .A1(n145), .A2(ctrl_DIV), .B1(n896), .B2(
        \product_reg/memory_26__dff/n5 ), .ZN(n299) );
  NAND4_X2 U294 ( .A1(n131), .A2(n132), .A3(n418), .A4(n419), .ZN(n288) );
  NOR4_X2 U295 ( .A1(n404), .A2(n401), .A3(n402), .A4(n400), .ZN(n419) );
  AOI22_X2 U300 ( .A1(n161), .A2(ctrl_DIV), .B1(n896), .B2(
        \product_reg/memory_10__dff/n5 ), .ZN(n339) );
  NAND2_X2 U301 ( .A1(n341), .A2(n340), .ZN(n338) );
  OAI22_X2 U302 ( .A1(data_operandA[8]), .A2(n896), .B1(ctrl_DIV), .B2(
        product_out[9]), .ZN(n340) );
  AOI22_X2 U304 ( .A1(n163), .A2(ctrl_DIV), .B1(n896), .B2(
        \product_reg/memory_8__dff/n5 ), .ZN(n343) );
  AOI22_X2 U307 ( .A1(n166), .A2(ctrl_DIV), .B1(n896), .B2(
        \product_reg/memory_5__dff/n5 ), .ZN(n320) );
  NAND2_X2 U308 ( .A1(n323), .A2(n122), .ZN(n319) );
  AOI22_X2 U309 ( .A1(n167), .A2(ctrl_DIV), .B1(n896), .B2(
        \product_reg/memory_4__dff/n5 ), .ZN(n322) );
  AOI22_X2 U311 ( .A1(n168), .A2(ctrl_DIV), .B1(n896), .B2(
        \product_reg/memory_3__dff/n5 ), .ZN(n317) );
  NAND2_X2 U312 ( .A1(n325), .A2(n326), .ZN(n316) );
  AOI22_X2 U313 ( .A1(ctrl_DIV), .A2(data_operandA[1]), .B1(product_out[2]), 
        .B2(n895), .ZN(n326) );
  AOI22_X2 U314 ( .A1(ctrl_DIV), .A2(data_operandA[0]), .B1(n120), .B2(n895), 
        .ZN(n325) );
  OAI22_X2 U315 ( .A1(data_operandA[5]), .A2(n896), .B1(ctrl_DIV), .B2(
        product_out[6]), .ZN(n346) );
  AOI22_X2 U316 ( .A1(n164), .A2(ctrl_DIV), .B1(n896), .B2(
        \product_reg/memory_7__dff/n5 ), .ZN(n420) );
  AOI22_X2 U317 ( .A1(n159), .A2(ctrl_DIV), .B1(n896), .B2(
        \product_reg/memory_12__dff/n5 ), .ZN(n421) );
  AOI22_X2 U318 ( .A1(n160), .A2(ctrl_DIV), .B1(n896), .B2(
        \product_reg/memory_11__dff/n5 ), .ZN(n415) );
  AOI22_X2 U319 ( .A1(n158), .A2(ctrl_DIV), .B1(n896), .B2(
        \product_reg/memory_13__dff/n5 ), .ZN(n410) );
  AOI22_X2 U320 ( .A1(n157), .A2(ctrl_DIV), .B1(n896), .B2(
        \product_reg/memory_14__dff/n5 ), .ZN(n408) );
  AOI22_X2 U321 ( .A1(n156), .A2(ctrl_DIV), .B1(n895), .B2(
        \product_reg/memory_15__dff/n5 ), .ZN(n412) );
  AOI22_X2 U322 ( .A1(n155), .A2(ctrl_DIV), .B1(n895), .B2(
        \product_reg/memory_16__dff/n5 ), .ZN(n422) );
  AOI22_X2 U323 ( .A1(n153), .A2(ctrl_DIV), .B1(n895), .B2(
        \product_reg/memory_18__dff/n5 ), .ZN(n402) );
  AOI22_X2 U324 ( .A1(n154), .A2(ctrl_DIV), .B1(n896), .B2(
        \product_reg/memory_17__dff/n5 ), .ZN(n401) );
  AOI22_X2 U325 ( .A1(n152), .A2(ctrl_DIV), .B1(n895), .B2(
        \product_reg/memory_19__dff/n5 ), .ZN(n404) );
  AOI22_X2 U327 ( .A1(n148), .A2(ctrl_DIV), .B1(n895), .B2(
        \product_reg/memory_23__dff/n5 ), .ZN(n304) );
  AOI22_X2 U328 ( .A1(n147), .A2(ctrl_DIV), .B1(n895), .B2(
        \product_reg/memory_24__dff/n5 ), .ZN(n302) );
  AOI22_X2 U329 ( .A1(n150), .A2(ctrl_DIV), .B1(n895), .B2(
        \product_reg/memory_21__dff/n5 ), .ZN(n348) );
  AOI22_X2 U330 ( .A1(n149), .A2(ctrl_DIV), .B1(n895), .B2(
        \product_reg/memory_22__dff/n5 ), .ZN(n347) );
  AOI22_X2 U331 ( .A1(n151), .A2(ctrl_DIV), .B1(n895), .B2(
        \product_reg/memory_20__dff/n5 ), .ZN(n423) );
  AOI22_X2 U332 ( .A1(n146), .A2(ctrl_DIV), .B1(n895), .B2(
        \product_reg/memory_25__dff/n5 ), .ZN(n289) );
  AOI22_X2 U333 ( .A1(n144), .A2(ctrl_DIV), .B1(n895), .B2(
        \product_reg/memory_27__dff/n5 ), .ZN(n292) );
  AOI22_X2 U334 ( .A1(n143), .A2(ctrl_DIV), .B1(n895), .B2(
        \product_reg/memory_28__dff/n5 ), .ZN(n296) );
  AOI22_X2 U335 ( .A1(n141), .A2(ctrl_DIV), .B1(n895), .B2(
        \product_reg/memory_30__dff/n5 ), .ZN(n283) );
  AOI22_X2 U336 ( .A1(n142), .A2(ctrl_DIV), .B1(n895), .B2(
        \product_reg/memory_29__dff/n5 ), .ZN(n285) );
  XNOR2_X2 U338 ( .A(n171), .B(data_operandA[31]), .ZN(n366) );
  NAND2_X2 U341 ( .A1(n758), .A2(n878), .ZN(n424) );
  OAI22_X2 U342 ( .A1(n845), .A2(\ctrl/mult_ready ), .B1(n850), .B2(n762), 
        .ZN(n216) );
  XNOR2_X2 U343 ( .A(n425), .B(n426), .ZN(adder_out[9]) );
  OAI22_X2 U345 ( .A1(n429), .A2(n430), .B1(n78), .B2(n431), .ZN(adder_out[8])
         );
  XNOR2_X2 U346 ( .A(n432), .B(n433), .ZN(n431) );
  XNOR2_X2 U348 ( .A(n436), .B(n437), .ZN(adder_out[7]) );
  XNOR2_X2 U349 ( .A(n438), .B(n439), .ZN(n437) );
  XOR2_X2 U350 ( .A(n440), .B(n441), .Z(adder_out[6]) );
  NAND2_X2 U351 ( .A1(n86), .A2(n442), .ZN(n440) );
  XNOR2_X2 U354 ( .A(n449), .B(n450), .ZN(n445) );
  OAI22_X2 U355 ( .A1(n451), .A2(n452), .B1(n80), .B2(n453), .ZN(adder_out[4])
         );
  XNOR2_X2 U356 ( .A(n454), .B(n455), .ZN(n453) );
  XNOR2_X2 U358 ( .A(n457), .B(n458), .ZN(adder_out[3]) );
  XNOR2_X2 U359 ( .A(n459), .B(n460), .ZN(n458) );
  XOR2_X2 U360 ( .A(n461), .B(n462), .Z(n748) );
  XOR2_X2 U362 ( .A(n466), .B(n467), .Z(n461) );
  OAI22_X2 U363 ( .A1(n850), .A2(\product_reg/memory_63__dff/n6 ), .B1(n847), 
        .B2(\product_reg/memory_64__dff/n5 ), .ZN(n467) );
  AOI221_X2 U364 ( .B1(n468), .B2(n469), .C1(n470), .C2(n864), .A(n887), .ZN(
        n466) );
  OAI221_X2 U365 ( .B1(n862), .B2(n171), .C1(n859), .C2(n897), .A(n473), .ZN(
        n469) );
  AOI22_X2 U366 ( .A1(n897), .A2(n854), .B1(n171), .B2(n853), .ZN(n473) );
  XOR2_X2 U367 ( .A(n463), .B(n476), .Z(adder_out[30]) );
  AND2_X2 U369 ( .A1(n477), .A2(n478), .ZN(n464) );
  AOI221_X2 U371 ( .B1(n866), .B2(n470), .C1(n479), .C2(n863), .A(n887), .ZN(
        n477) );
  OAI221_X2 U372 ( .B1(n862), .B2(n172), .C1(n859), .C2(n140), .A(n480), .ZN(
        n470) );
  AOI22_X2 U373 ( .A1(n853), .A2(n172), .B1(n854), .B2(n140), .ZN(n480) );
  AOI22_X2 U374 ( .A1(n849), .A2(\product_reg/memory_63__dff/n6 ), .B1(n846), 
        .B2(\product_reg/memory_62__dff/n5 ), .ZN(n478) );
  OAI22_X2 U377 ( .A1(n485), .A2(n486), .B1(n81), .B2(n487), .ZN(adder_out[2])
         );
  XNOR2_X2 U378 ( .A(n488), .B(n489), .ZN(n487) );
  OAI221_X2 U380 ( .B1(n484), .B2(n492), .C1(n72), .C2(n482), .A(n493), .ZN(
        adder_out[29]) );
  NAND2_X2 U382 ( .A1(n483), .A2(n484), .ZN(n482) );
  XOR2_X2 U383 ( .A(n72), .B(n483), .Z(n492) );
  AOI221_X2 U384 ( .B1(n468), .B2(n479), .C1(n494), .C2(n863), .A(n887), .ZN(
        n483) );
  OAI221_X2 U385 ( .B1(n862), .B2(n173), .C1(n141), .C2(n857), .A(n495), .ZN(
        n479) );
  AOI22_X2 U386 ( .A1(n853), .A2(n173), .B1(n854), .B2(n141), .ZN(n495) );
  OAI22_X2 U389 ( .A1(\product_reg/memory_62__dff/n5 ), .A2(n847), .B1(
        \product_reg/memory_61__dff/n5 ), .B2(n850), .ZN(n484) );
  OAI221_X2 U390 ( .B1(n500), .B2(n501), .C1(n73), .C2(n498), .A(n502), .ZN(
        adder_out[28]) );
  NAND2_X2 U392 ( .A1(n499), .A2(n500), .ZN(n498) );
  XOR2_X2 U393 ( .A(n107), .B(n503), .Z(n501) );
  AOI221_X2 U395 ( .B1(n468), .B2(n494), .C1(n507), .C2(n863), .A(n887), .ZN(
        n499) );
  OAI221_X2 U396 ( .B1(n862), .B2(n174), .C1(n142), .C2(n857), .A(n508), .ZN(
        n494) );
  AOI22_X2 U397 ( .A1(n853), .A2(n174), .B1(n854), .B2(n142), .ZN(n508) );
  OAI22_X2 U398 ( .A1(\product_reg/memory_61__dff/n5 ), .A2(n847), .B1(
        \product_reg/memory_60__dff/n5 ), .B2(n850), .ZN(n500) );
  XOR2_X2 U399 ( .A(n509), .B(n504), .Z(adder_out[27]) );
  NAND2_X2 U401 ( .A1(n105), .A2(n112), .ZN(n510) );
  NAND2_X2 U402 ( .A1(n506), .A2(n106), .ZN(n509) );
  NAND2_X2 U404 ( .A1(n513), .A2(n512), .ZN(n506) );
  AOI22_X2 U405 ( .A1(n849), .A2(\product_reg/memory_60__dff/n5 ), .B1(n845), 
        .B2(\product_reg/memory_59__dff/n5 ), .ZN(n512) );
  AOI221_X2 U406 ( .B1(n468), .B2(n507), .C1(n514), .C2(n863), .A(n887), .ZN(
        n513) );
  OAI221_X2 U407 ( .B1(n862), .B2(n175), .C1(n143), .C2(n857), .A(n515), .ZN(
        n507) );
  AOI22_X2 U408 ( .A1(n853), .A2(n175), .B1(n854), .B2(n143), .ZN(n515) );
  OAI22_X2 U409 ( .A1(n516), .A2(n517), .B1(n74), .B2(n518), .ZN(adder_out[26]) );
  XOR2_X2 U410 ( .A(n105), .B(n519), .Z(n518) );
  AOI221_X2 U413 ( .B1(n468), .B2(n514), .C1(n521), .C2(n863), .A(n887), .ZN(
        n520) );
  OAI221_X2 U414 ( .B1(n862), .B2(n176), .C1(n144), .C2(n857), .A(n522), .ZN(
        n514) );
  AOI22_X2 U415 ( .A1(n853), .A2(n176), .B1(n854), .B2(n144), .ZN(n522) );
  OAI22_X2 U416 ( .A1(\product_reg/memory_59__dff/n5 ), .A2(n847), .B1(
        \product_reg/memory_58__dff/n5 ), .B2(n850), .ZN(n519) );
  XOR2_X2 U418 ( .A(n523), .B(n526), .Z(adder_out[25]) );
  AND2_X2 U420 ( .A1(n527), .A2(n528), .ZN(n524) );
  AOI221_X2 U422 ( .B1(n468), .B2(n521), .C1(n529), .C2(n863), .A(n887), .ZN(
        n527) );
  OAI221_X2 U423 ( .B1(n862), .B2(n177), .C1(n145), .C2(n857), .A(n530), .ZN(
        n521) );
  AOI22_X2 U424 ( .A1(n853), .A2(n177), .B1(n854), .B2(n145), .ZN(n530) );
  AOI22_X2 U425 ( .A1(n849), .A2(\product_reg/memory_58__dff/n5 ), .B1(n845), 
        .B2(\product_reg/memory_57__dff/n5 ), .ZN(n528) );
  OAI221_X2 U428 ( .B1(n535), .B2(n536), .C1(n532), .C2(n533), .A(n537), .ZN(
        adder_out[24]) );
  NAND2_X2 U430 ( .A1(n534), .A2(n535), .ZN(n533) );
  XOR2_X2 U431 ( .A(n534), .B(n532), .Z(n536) );
  AOI22_X2 U432 ( .A1(n538), .A2(n539), .B1(n102), .B2(n540), .ZN(n532) );
  AOI221_X2 U433 ( .B1(n468), .B2(n529), .C1(n542), .C2(n864), .A(n887), .ZN(
        n534) );
  OAI221_X2 U434 ( .B1(n862), .B2(n178), .C1(n146), .C2(n857), .A(n543), .ZN(
        n529) );
  AOI22_X2 U435 ( .A1(n853), .A2(n178), .B1(n854), .B2(n146), .ZN(n543) );
  OAI22_X2 U436 ( .A1(\product_reg/memory_57__dff/n5 ), .A2(n846), .B1(
        \product_reg/memory_56__dff/n5 ), .B2(n850), .ZN(n535) );
  XOR2_X2 U437 ( .A(n540), .B(n544), .Z(adder_out[23]) );
  OAI22_X2 U440 ( .A1(\product_reg/memory_56__dff/n5 ), .A2(n846), .B1(
        \product_reg/memory_55__dff/n5 ), .B2(n850), .ZN(n538) );
  AOI221_X2 U441 ( .B1(n468), .B2(n542), .C1(n545), .C2(n864), .A(n887), .ZN(
        n539) );
  OAI221_X2 U442 ( .B1(n862), .B2(n179), .C1(n147), .C2(n858), .A(n546), .ZN(
        n542) );
  AOI22_X2 U443 ( .A1(n853), .A2(n179), .B1(n854), .B2(n147), .ZN(n546) );
  XNOR2_X2 U445 ( .A(n548), .B(n550), .ZN(adder_out[22]) );
  NAND2_X2 U447 ( .A1(n551), .A2(n552), .ZN(n549) );
  AOI221_X2 U449 ( .B1(n468), .B2(n545), .C1(n553), .C2(n864), .A(n887), .ZN(
        n551) );
  OAI221_X2 U450 ( .B1(n862), .B2(n180), .C1(n859), .C2(n148), .A(n554), .ZN(
        n545) );
  AOI22_X2 U451 ( .A1(n853), .A2(n180), .B1(n854), .B2(n148), .ZN(n554) );
  AOI22_X2 U452 ( .A1(n849), .A2(\product_reg/memory_55__dff/n5 ), .B1(n845), 
        .B2(\product_reg/memory_54__dff/n5 ), .ZN(n552) );
  XOR2_X2 U454 ( .A(n555), .B(n558), .Z(adder_out[21]) );
  AND2_X2 U456 ( .A1(n559), .A2(n560), .ZN(n556) );
  AOI221_X2 U458 ( .B1(n468), .B2(n553), .C1(n561), .C2(n864), .A(n887), .ZN(
        n559) );
  OAI221_X2 U459 ( .B1(n861), .B2(n181), .C1(n858), .C2(n149), .A(n562), .ZN(
        n553) );
  AOI22_X2 U460 ( .A1(n852), .A2(n181), .B1(n854), .B2(n149), .ZN(n562) );
  OAI22_X2 U461 ( .A1(\product_reg/memory_54__dff/n5 ), .A2(n846), .B1(
        \product_reg/memory_53__dff/n5 ), .B2(n850), .ZN(n560) );
  OAI22_X2 U463 ( .A1(n75), .A2(n565), .B1(n566), .B2(n567), .ZN(adder_out[20]) );
  XNOR2_X2 U464 ( .A(n568), .B(n569), .ZN(n567) );
  NAND2_X2 U466 ( .A1(n569), .A2(n568), .ZN(n564) );
  AOI221_X2 U468 ( .B1(n866), .B2(n561), .C1(n570), .C2(n864), .A(n888), .ZN(
        n569) );
  OAI221_X2 U469 ( .B1(n861), .B2(n182), .C1(n857), .C2(n150), .A(n571), .ZN(
        n561) );
  AOI22_X2 U470 ( .A1(n852), .A2(n182), .B1(n855), .B2(n150), .ZN(n571) );
  OAI22_X2 U471 ( .A1(\product_reg/memory_53__dff/n5 ), .A2(n846), .B1(
        \product_reg/memory_52__dff/n5 ), .B2(n850), .ZN(n568) );
  XOR2_X2 U473 ( .A(n113), .B(n575), .Z(adder_out[1]) );
  XOR2_X2 U474 ( .A(n576), .B(n577), .Z(n575) );
  XNOR2_X2 U475 ( .A(n572), .B(n578), .ZN(adder_out[19]) );
  NAND2_X2 U477 ( .A1(n579), .A2(n580), .ZN(n574) );
  AOI221_X2 U479 ( .B1(n867), .B2(n570), .C1(n581), .C2(n864), .A(n888), .ZN(
        n579) );
  OAI221_X2 U480 ( .B1(n861), .B2(n183), .C1(n151), .C2(n857), .A(n582), .ZN(
        n570) );
  AOI22_X2 U481 ( .A1(n852), .A2(n183), .B1(n855), .B2(n151), .ZN(n582) );
  AOI22_X2 U482 ( .A1(n849), .A2(\product_reg/memory_52__dff/n5 ), .B1(n845), 
        .B2(\product_reg/memory_51__dff/n5 ), .ZN(n580) );
  OAI22_X2 U484 ( .A1(n585), .A2(n586), .B1(n76), .B2(n587), .ZN(adder_out[18]) );
  XNOR2_X2 U485 ( .A(n588), .B(n589), .ZN(n587) );
  AND2_X2 U487 ( .A1(n588), .A2(n589), .ZN(n583) );
  AOI221_X2 U489 ( .B1(n867), .B2(n581), .C1(n590), .C2(n864), .A(n888), .ZN(
        n588) );
  OAI221_X2 U490 ( .B1(n861), .B2(n184), .C1(n152), .C2(n857), .A(n591), .ZN(
        n581) );
  AOI22_X2 U491 ( .A1(n852), .A2(n184), .B1(n855), .B2(n152), .ZN(n591) );
  OAI22_X2 U492 ( .A1(\product_reg/memory_51__dff/n5 ), .A2(n846), .B1(
        \product_reg/memory_50__dff/n5 ), .B2(n850), .ZN(n589) );
  XOR2_X2 U494 ( .A(n592), .B(n595), .Z(adder_out[17]) );
  AND2_X2 U496 ( .A1(n596), .A2(n597), .ZN(n593) );
  AOI221_X2 U498 ( .B1(n867), .B2(n590), .C1(n598), .C2(n864), .A(n888), .ZN(
        n596) );
  OAI221_X2 U499 ( .B1(n861), .B2(n185), .C1(n153), .C2(n857), .A(n599), .ZN(
        n590) );
  AOI22_X2 U500 ( .A1(n852), .A2(n185), .B1(n855), .B2(n153), .ZN(n599) );
  AOI22_X2 U501 ( .A1(n849), .A2(\product_reg/memory_50__dff/n5 ), .B1(n845), 
        .B2(\product_reg/memory_49__dff/n5 ), .ZN(n597) );
  OAI22_X2 U503 ( .A1(n601), .A2(n603), .B1(n70), .B2(n604), .ZN(adder_out[16]) );
  XNOR2_X2 U504 ( .A(n605), .B(n606), .ZN(n604) );
  NAND2_X2 U506 ( .A1(n606), .A2(n605), .ZN(n602) );
  AOI221_X2 U508 ( .B1(n867), .B2(n598), .C1(n607), .C2(n864), .A(n888), .ZN(
        n606) );
  OAI221_X2 U509 ( .B1(n861), .B2(n186), .C1(n154), .C2(n857), .A(n608), .ZN(
        n598) );
  AOI22_X2 U510 ( .A1(n852), .A2(n186), .B1(n855), .B2(n154), .ZN(n608) );
  OAI22_X2 U511 ( .A1(\product_reg/memory_49__dff/n5 ), .A2(n846), .B1(
        \product_reg/memory_48__dff/n5 ), .B2(n850), .ZN(n605) );
  AOI22_X2 U512 ( .A1(n609), .A2(n610), .B1(n94), .B2(n611), .ZN(n601) );
  XOR2_X2 U513 ( .A(n611), .B(n613), .Z(adder_out[15]) );
  OAI22_X2 U516 ( .A1(\product_reg/memory_48__dff/n5 ), .A2(n846), .B1(
        \product_reg/memory_47__dff/n5 ), .B2(n850), .ZN(n609) );
  AOI221_X2 U517 ( .B1(n867), .B2(n607), .C1(n614), .C2(n863), .A(n888), .ZN(
        n610) );
  OAI221_X2 U518 ( .B1(n861), .B2(n188), .C1(n155), .C2(n858), .A(n615), .ZN(
        n607) );
  AOI22_X2 U519 ( .A1(n852), .A2(n188), .B1(n855), .B2(n155), .ZN(n615) );
  XNOR2_X2 U521 ( .A(n617), .B(n619), .ZN(adder_out[14]) );
  NAND2_X2 U523 ( .A1(n620), .A2(n621), .ZN(n618) );
  AOI221_X2 U525 ( .B1(n867), .B2(n614), .C1(n622), .C2(n863), .A(n888), .ZN(
        n620) );
  OAI221_X2 U526 ( .B1(n861), .B2(n189), .C1(n156), .C2(n858), .A(n623), .ZN(
        n614) );
  AOI22_X2 U527 ( .A1(n852), .A2(n189), .B1(n855), .B2(n156), .ZN(n623) );
  AOI22_X2 U528 ( .A1(n849), .A2(\product_reg/memory_47__dff/n5 ), .B1(n845), 
        .B2(\product_reg/memory_46__dff/n5 ), .ZN(n621) );
  XOR2_X2 U530 ( .A(n624), .B(n628), .Z(adder_out[13]) );
  AND2_X2 U532 ( .A1(n629), .A2(n630), .ZN(n626) );
  AOI221_X2 U534 ( .B1(n867), .B2(n622), .C1(n631), .C2(n863), .A(n888), .ZN(
        n629) );
  OAI221_X2 U535 ( .B1(n861), .B2(n190), .C1(n157), .C2(n858), .A(n632), .ZN(
        n622) );
  AOI22_X2 U536 ( .A1(n852), .A2(n190), .B1(n855), .B2(n157), .ZN(n632) );
  OAI22_X2 U537 ( .A1(\product_reg/memory_46__dff/n5 ), .A2(n846), .B1(
        \product_reg/memory_45__dff/n5 ), .B2(n850), .ZN(n630) );
  OAI22_X2 U539 ( .A1(n77), .A2(n635), .B1(n636), .B2(n637), .ZN(adder_out[12]) );
  XNOR2_X2 U540 ( .A(n638), .B(n639), .ZN(n637) );
  NAND2_X2 U542 ( .A1(n639), .A2(n638), .ZN(n634) );
  AOI221_X2 U544 ( .B1(n867), .B2(n631), .C1(n640), .C2(n863), .A(n888), .ZN(
        n639) );
  OAI221_X2 U545 ( .B1(n861), .B2(n191), .C1(n158), .C2(n858), .A(n641), .ZN(
        n631) );
  AOI22_X2 U546 ( .A1(n852), .A2(n191), .B1(n855), .B2(n158), .ZN(n641) );
  OAI22_X2 U547 ( .A1(\product_reg/memory_45__dff/n5 ), .A2(n846), .B1(
        \product_reg/memory_44__dff/n5 ), .B2(n849), .ZN(n638) );
  XNOR2_X2 U549 ( .A(n642), .B(n645), .ZN(adder_out[11]) );
  NAND2_X2 U551 ( .A1(n646), .A2(n647), .ZN(n644) );
  AOI221_X2 U553 ( .B1(n867), .B2(n640), .C1(n648), .C2(n865), .A(n888), .ZN(
        n646) );
  OAI221_X2 U554 ( .B1(n861), .B2(n192), .C1(n159), .C2(n858), .A(n649), .ZN(
        n640) );
  AOI22_X2 U555 ( .A1(n852), .A2(n192), .B1(n855), .B2(n159), .ZN(n649) );
  AOI22_X2 U556 ( .A1(n849), .A2(\product_reg/memory_44__dff/n5 ), .B1(n845), 
        .B2(\product_reg/memory_43__dff/n5 ), .ZN(n647) );
  OAI22_X2 U558 ( .A1(n69), .A2(n653), .B1(n650), .B2(n654), .ZN(adder_out[10]) );
  XNOR2_X2 U559 ( .A(n655), .B(n656), .ZN(n654) );
  AND2_X2 U561 ( .A1(n655), .A2(n656), .ZN(n651) );
  AOI221_X2 U563 ( .B1(n867), .B2(n648), .C1(n657), .C2(n865), .A(n888), .ZN(
        n655) );
  OAI221_X2 U564 ( .B1(n860), .B2(n193), .C1(n160), .C2(n858), .A(n658), .ZN(
        n648) );
  AOI22_X2 U565 ( .A1(n851), .A2(n193), .B1(n855), .B2(n160), .ZN(n658) );
  OAI22_X2 U566 ( .A1(\product_reg/memory_43__dff/n5 ), .A2(n846), .B1(
        \product_reg/memory_42__dff/n5 ), .B2(n849), .ZN(n656) );
  NAND2_X2 U568 ( .A1(n659), .A2(n660), .ZN(n428) );
  AND2_X2 U570 ( .A1(n432), .A2(n433), .ZN(n435) );
  NAND2_X2 U574 ( .A1(n662), .A2(n663), .ZN(n442) );
  AND2_X2 U576 ( .A1(n449), .A2(n450), .ZN(n448) );
  AOI22_X2 U579 ( .A1(n459), .A2(n457), .B1(n665), .B2(n460), .ZN(n451) );
  NAND2_X2 U581 ( .A1(n488), .A2(n489), .ZN(n491) );
  NAND2_X2 U584 ( .A1(n668), .A2(n669), .ZN(n576) );
  OAI22_X2 U585 ( .A1(n867), .A2(n670), .B1(n865), .B2(n671), .ZN(n668) );
  OAI22_X2 U586 ( .A1(\product_reg/memory_34__dff/n5 ), .A2(n846), .B1(
        \product_reg/memory_33__dff/n5 ), .B2(n850), .ZN(n666) );
  AOI221_X2 U589 ( .B1(n867), .B2(n674), .C1(n671), .C2(n863), .A(n889), .ZN(
        n488) );
  OAI221_X2 U590 ( .B1(n860), .B2(n205), .C1(n169), .C2(n858), .A(n675), .ZN(
        n671) );
  AOI22_X2 U591 ( .A1(n851), .A2(n205), .B1(n856), .B2(n169), .ZN(n675) );
  OAI22_X2 U592 ( .A1(\product_reg/memory_35__dff/n5 ), .A2(n846), .B1(
        \product_reg/memory_34__dff/n5 ), .B2(n849), .ZN(n489) );
  OR2_X2 U593 ( .A1(n457), .A2(n459), .ZN(n665) );
  AOI221_X2 U594 ( .B1(n867), .B2(n676), .C1(n674), .C2(n865), .A(n889), .ZN(
        n457) );
  OAI221_X2 U595 ( .B1(n860), .B2(n204), .C1(n168), .C2(n858), .A(n677), .ZN(
        n674) );
  AOI22_X2 U596 ( .A1(n851), .A2(n204), .B1(n856), .B2(n168), .ZN(n677) );
  OAI22_X2 U597 ( .A1(\product_reg/memory_36__dff/n5 ), .A2(n846), .B1(
        \product_reg/memory_35__dff/n5 ), .B2(n850), .ZN(n459) );
  NAND2_X2 U598 ( .A1(n455), .A2(n454), .ZN(n664) );
  AOI221_X2 U599 ( .B1(n867), .B2(n678), .C1(n676), .C2(n865), .A(n889), .ZN(
        n454) );
  OAI221_X2 U600 ( .B1(n860), .B2(n203), .C1(n167), .C2(n858), .A(n679), .ZN(
        n676) );
  AOI22_X2 U601 ( .A1(n851), .A2(n203), .B1(n856), .B2(n167), .ZN(n679) );
  OAI22_X2 U602 ( .A1(\product_reg/memory_37__dff/n5 ), .A2(n846), .B1(
        \product_reg/memory_36__dff/n5 ), .B2(n850), .ZN(n455) );
  AOI221_X2 U604 ( .B1(n867), .B2(n680), .C1(n678), .C2(n865), .A(n889), .ZN(
        n449) );
  OAI221_X2 U605 ( .B1(n860), .B2(n202), .C1(n166), .C2(n858), .A(n681), .ZN(
        n678) );
  AOI22_X2 U606 ( .A1(n851), .A2(n202), .B1(n856), .B2(n166), .ZN(n681) );
  OAI22_X2 U607 ( .A1(\product_reg/memory_38__dff/n5 ), .A2(n846), .B1(
        \product_reg/memory_37__dff/n5 ), .B2(n849), .ZN(n450) );
  AOI221_X2 U609 ( .B1(n867), .B2(n682), .C1(n680), .C2(n865), .A(n889), .ZN(
        n662) );
  OAI221_X2 U610 ( .B1(n860), .B2(n201), .C1(n859), .C2(n165), .A(n683), .ZN(
        n680) );
  AOI22_X2 U611 ( .A1(n851), .A2(n201), .B1(n856), .B2(n165), .ZN(n683) );
  AOI22_X2 U612 ( .A1(n849), .A2(\product_reg/memory_39__dff/n5 ), .B1(n845), 
        .B2(\product_reg/memory_38__dff/n5 ), .ZN(n663) );
  AOI221_X2 U613 ( .B1(n867), .B2(n684), .C1(n682), .C2(n864), .A(n889), .ZN(
        n439) );
  OAI221_X2 U614 ( .B1(n860), .B2(n200), .C1(n859), .C2(n164), .A(n685), .ZN(
        n682) );
  AOI22_X2 U615 ( .A1(n851), .A2(n200), .B1(n856), .B2(n164), .ZN(n685) );
  OAI22_X2 U616 ( .A1(\product_reg/memory_40__dff/n5 ), .A2(n847), .B1(
        \product_reg/memory_39__dff/n5 ), .B2(n849), .ZN(n436) );
  AOI221_X2 U618 ( .B1(n867), .B2(n686), .C1(n684), .C2(n865), .A(n889), .ZN(
        n432) );
  OAI221_X2 U619 ( .B1(n860), .B2(n199), .C1(n859), .C2(n163), .A(n687), .ZN(
        n684) );
  AOI22_X2 U620 ( .A1(n851), .A2(n199), .B1(n856), .B2(n163), .ZN(n687) );
  OAI22_X2 U621 ( .A1(\product_reg/memory_41__dff/n5 ), .A2(n846), .B1(
        \product_reg/memory_40__dff/n5 ), .B2(n849), .ZN(n433) );
  AOI221_X2 U623 ( .B1(n867), .B2(n657), .C1(n686), .C2(n864), .A(n889), .ZN(
        n659) );
  OAI221_X2 U624 ( .B1(n860), .B2(n195), .C1(n859), .C2(n162), .A(n688), .ZN(
        n686) );
  AOI22_X2 U625 ( .A1(n851), .A2(n195), .B1(n856), .B2(n162), .ZN(n688) );
  OAI221_X2 U626 ( .B1(n860), .B2(n194), .C1(n859), .C2(n161), .A(n689), .ZN(
        n657) );
  AOI22_X2 U627 ( .A1(n851), .A2(n194), .B1(n856), .B2(n161), .ZN(n689) );
  AOI22_X2 U628 ( .A1(n848), .A2(\product_reg/memory_42__dff/n5 ), .B1(n845), 
        .B2(\product_reg/memory_41__dff/n5 ), .ZN(n660) );
  OAI22_X2 U629 ( .A1(n115), .A2(n690), .B1(n691), .B2(n692), .ZN(adder_out[0]) );
  XNOR2_X2 U630 ( .A(n693), .B(n694), .ZN(n692) );
  NAND2_X2 U632 ( .A1(n694), .A2(n693), .ZN(n673) );
  AOI221_X2 U634 ( .B1(n115), .B2(n863), .C1(n867), .C2(n670), .A(n889), .ZN(
        n694) );
  NAND4_X2 U635 ( .A1(\ctrl/op_mult_int ), .A2(n695), .A3(n696), .A4(n697), 
        .ZN(n669) );
  OAI221_X2 U637 ( .B1(n860), .B2(n206), .C1(n170), .C2(n857), .A(n698), .ZN(
        n670) );
  AOI22_X2 U638 ( .A1(n851), .A2(n206), .B1(n856), .B2(n170), .ZN(n698) );
  NAND2_X2 U643 ( .A1(\ctrl/op_mult_int ), .A2(n699), .ZN(n468) );
  NAND2_X2 U646 ( .A1(\product_reg/memory_2__dff/n7 ), .A2(n120), .ZN(n697) );
  OAI22_X2 U647 ( .A1(\product_reg/memory_33__dff/n5 ), .A2(n846), .B1(n850), 
        .B2(n135), .ZN(n693) );
  OAI22_X2 U650 ( .A1(\ctrl/op_mult_int ), .A2(n701), .B1(n695), .B2(n116), 
        .ZN(n691) );
  XOR2_X2 U652 ( .A(n171), .B(\product_reg/memory_63__dff/n6 ), .Z(n701) );
  INV_X4 U653 ( .A(n279), .ZN(n65) );
  INV_X4 U657 ( .A(n650), .ZN(n69) );
  INV_X4 U658 ( .A(n601), .ZN(n70) );
  INV_X4 U659 ( .A(n748), .ZN(n71) );
  INV_X4 U660 ( .A(n496), .ZN(n72) );
  INV_X4 U661 ( .A(n503), .ZN(n73) );
  INV_X4 U662 ( .A(n516), .ZN(n74) );
  INV_X4 U663 ( .A(n566), .ZN(n75) );
  INV_X4 U664 ( .A(n585), .ZN(n76) );
  INV_X4 U665 ( .A(n636), .ZN(n77) );
  INV_X4 U666 ( .A(n429), .ZN(n78) );
  INV_X4 U667 ( .A(n661), .ZN(n79) );
  INV_X4 U668 ( .A(n451), .ZN(n80) );
  INV_X4 U669 ( .A(n485), .ZN(n81) );
  INV_X4 U670 ( .A(n577), .ZN(n82) );
  INV_X4 U671 ( .A(n673), .ZN(n83) );
  INV_X4 U672 ( .A(n428), .ZN(n84) );
  INV_X4 U673 ( .A(n434), .ZN(n85) );
  INV_X4 U674 ( .A(n443), .ZN(n86) );
  INV_X4 U675 ( .A(n447), .ZN(n87) );
  INV_X4 U676 ( .A(n491), .ZN(n88) );
  INV_X4 U677 ( .A(n652), .ZN(n89) );
  INV_X4 U678 ( .A(n644), .ZN(n90) );
  INV_X4 U679 ( .A(n634), .ZN(n91) );
  INV_X4 U680 ( .A(n627), .ZN(n92) );
  INV_X4 U681 ( .A(n618), .ZN(n93) );
  INV_X4 U682 ( .A(n612), .ZN(n94) );
  INV_X4 U683 ( .A(n602), .ZN(n95) );
  INV_X4 U684 ( .A(n594), .ZN(n96) );
  INV_X4 U685 ( .A(n584), .ZN(n97) );
  INV_X4 U686 ( .A(n574), .ZN(n98) );
  INV_X4 U687 ( .A(n564), .ZN(n99) );
  INV_X4 U688 ( .A(n557), .ZN(n100) );
  INV_X4 U689 ( .A(n549), .ZN(n101) );
  INV_X4 U690 ( .A(n541), .ZN(n102) );
  INV_X4 U691 ( .A(n534), .ZN(n103) );
  INV_X4 U692 ( .A(n525), .ZN(n104) );
  INV_X4 U693 ( .A(n520), .ZN(n105) );
  INV_X4 U694 ( .A(n505), .ZN(n106) );
  INV_X4 U695 ( .A(n499), .ZN(n107) );
  INV_X4 U696 ( .A(n483), .ZN(n108) );
  INV_X4 U697 ( .A(n465), .ZN(n109) );
  INV_X4 U700 ( .A(n519), .ZN(n112) );
  INV_X4 U701 ( .A(n666), .ZN(n113) );
  INV_X4 U703 ( .A(n691), .ZN(n115) );
  INV_X4 U707 ( .A(n416), .ZN(n119) );
  INV_X4 U710 ( .A(n322), .ZN(n122) );
  INV_X4 U712 ( .A(n420), .ZN(n124) );
  INV_X4 U714 ( .A(n415), .ZN(n126) );
  INV_X4 U715 ( .A(n421), .ZN(n127) );
  INV_X4 U716 ( .A(n412), .ZN(n128) );
  INV_X4 U717 ( .A(n422), .ZN(n129) );
  INV_X4 U718 ( .A(n404), .ZN(n130) );
  INV_X4 U719 ( .A(n423), .ZN(n131) );
  INV_X4 U720 ( .A(n347), .ZN(n132) );
  INV_X4 U721 ( .A(n304), .ZN(n133) );
  INV_X4 U726 ( .A(n366), .ZN(n138) );
  INV_X4 U728 ( .A(data_operandA[30]), .ZN(n140) );
  INV_X4 U729 ( .A(data_operandA[29]), .ZN(n141) );
  INV_X4 U730 ( .A(data_operandA[28]), .ZN(n142) );
  INV_X4 U731 ( .A(data_operandA[27]), .ZN(n143) );
  INV_X4 U732 ( .A(data_operandA[26]), .ZN(n144) );
  INV_X4 U733 ( .A(data_operandA[25]), .ZN(n145) );
  INV_X4 U734 ( .A(data_operandA[24]), .ZN(n146) );
  INV_X4 U735 ( .A(data_operandA[23]), .ZN(n147) );
  INV_X4 U736 ( .A(data_operandA[22]), .ZN(n148) );
  INV_X4 U737 ( .A(data_operandA[21]), .ZN(n149) );
  INV_X4 U738 ( .A(data_operandA[20]), .ZN(n150) );
  INV_X4 U739 ( .A(data_operandA[19]), .ZN(n151) );
  INV_X4 U740 ( .A(data_operandA[18]), .ZN(n152) );
  INV_X4 U741 ( .A(data_operandA[17]), .ZN(n153) );
  INV_X4 U742 ( .A(data_operandA[16]), .ZN(n154) );
  INV_X4 U743 ( .A(data_operandA[15]), .ZN(n155) );
  INV_X4 U744 ( .A(data_operandA[14]), .ZN(n156) );
  INV_X4 U745 ( .A(data_operandA[13]), .ZN(n157) );
  INV_X4 U746 ( .A(data_operandA[12]), .ZN(n158) );
  INV_X4 U747 ( .A(data_operandA[11]), .ZN(n159) );
  INV_X4 U748 ( .A(data_operandA[10]), .ZN(n160) );
  INV_X4 U749 ( .A(data_operandA[9]), .ZN(n161) );
  INV_X4 U750 ( .A(data_operandA[8]), .ZN(n162) );
  INV_X4 U751 ( .A(data_operandA[7]), .ZN(n163) );
  INV_X4 U752 ( .A(data_operandA[6]), .ZN(n164) );
  INV_X4 U753 ( .A(data_operandA[5]), .ZN(n165) );
  INV_X4 U754 ( .A(data_operandA[4]), .ZN(n166) );
  INV_X4 U755 ( .A(data_operandA[3]), .ZN(n167) );
  INV_X4 U756 ( .A(data_operandA[2]), .ZN(n168) );
  INV_X4 U757 ( .A(data_operandA[1]), .ZN(n169) );
  INV_X4 U758 ( .A(data_operandA[0]), .ZN(n170) );
  INV_X4 U759 ( .A(data_operandB[31]), .ZN(n171) );
  INV_X4 U760 ( .A(data_operandB[30]), .ZN(n172) );
  INV_X4 U761 ( .A(data_operandB[29]), .ZN(n173) );
  INV_X4 U762 ( .A(data_operandB[28]), .ZN(n174) );
  INV_X4 U763 ( .A(data_operandB[27]), .ZN(n175) );
  INV_X4 U764 ( .A(data_operandB[26]), .ZN(n176) );
  INV_X4 U765 ( .A(data_operandB[25]), .ZN(n177) );
  INV_X4 U766 ( .A(data_operandB[24]), .ZN(n178) );
  INV_X4 U767 ( .A(data_operandB[23]), .ZN(n179) );
  INV_X4 U768 ( .A(data_operandB[22]), .ZN(n180) );
  INV_X4 U769 ( .A(data_operandB[21]), .ZN(n181) );
  INV_X4 U770 ( .A(data_operandB[20]), .ZN(n182) );
  INV_X4 U771 ( .A(data_operandB[19]), .ZN(n183) );
  INV_X4 U772 ( .A(data_operandB[18]), .ZN(n184) );
  INV_X4 U773 ( .A(data_operandB[17]), .ZN(n185) );
  INV_X4 U774 ( .A(data_operandB[16]), .ZN(n186) );
  INV_X4 U775 ( .A(data_operandB[15]), .ZN(n188) );
  INV_X4 U776 ( .A(data_operandB[14]), .ZN(n189) );
  INV_X4 U777 ( .A(data_operandB[13]), .ZN(n190) );
  INV_X4 U778 ( .A(data_operandB[12]), .ZN(n191) );
  INV_X4 U779 ( .A(data_operandB[11]), .ZN(n192) );
  INV_X4 U780 ( .A(data_operandB[10]), .ZN(n193) );
  INV_X4 U781 ( .A(data_operandB[9]), .ZN(n194) );
  INV_X4 U782 ( .A(data_operandB[8]), .ZN(n195) );
  INV_X4 U783 ( .A(data_operandB[7]), .ZN(n199) );
  INV_X4 U784 ( .A(data_operandB[6]), .ZN(n200) );
  INV_X4 U785 ( .A(data_operandB[5]), .ZN(n201) );
  INV_X4 U786 ( .A(data_operandB[4]), .ZN(n202) );
  INV_X4 U787 ( .A(data_operandB[3]), .ZN(n203) );
  INV_X4 U788 ( .A(data_operandB[2]), .ZN(n204) );
  INV_X4 U789 ( .A(data_operandB[1]), .ZN(n205) );
  INV_X4 U790 ( .A(data_operandB[0]), .ZN(n206) );
  INV_X4 U791 ( .A(ctrl_MULT), .ZN(n207) );
  INV_X4 U793 ( .A(clock), .ZN(n211) );
  SDFFR_X2 \ctrl/counter/tff_0/dffe/q_reg  ( .D(n749), .SI(test_si1), .SE(
        test_se), .CK(n211), .RN(n758), .Q(test_so1), .QN(n749) );
  SDFFR_X2 \ctrl/counter/tff_1/dffe/q_reg  ( .D(n750), .SI(1'b0), .SE(1'b0), 
        .CK(n749), .RN(n758), .QN(n750) );
  SDFFR_X2 \ctrl/counter/tff_2/dffe/q_reg  ( .D(n751), .SI(1'b0), .SE(1'b0), 
        .CK(n750), .RN(n758), .QN(n751) );
  SDFFR_X2 \ctrl/counter/tff_3/dffe/q_reg  ( .D(n752), .SI(1'b0), .SE(1'b0), 
        .CK(n751), .RN(n758), .QN(n752) );
  SDFFR_X2 \ctrl/counter/tff_4/dffe/q_reg  ( .D(n753), .SI(1'b0), .SE(1'b0), 
        .CK(n752), .RN(n758), .Q(\ctrl/counter/w5 ), .QN(n753) );
  SDFFR_X2 \ctrl/counter/tff_5/dffe/q_reg  ( .D(n754), .SI(1'b0), .SE(1'b0), 
        .CK(n753), .RN(n758), .Q(\ctrl/counter/w7 ), .QN(n754) );
  SDFFR_X2 \ctrl/counter/output16_dff/q_reg  ( .D(\ctrl/counter/w5 ), .SI(
        test_si2), .SE(test_se), .CK(clock), .RN(n758), .Q(\ctrl/mult_ready ), 
        .QN(n1037) );
  SDFFR_X2 \ctrl/counter/output32_dff/q_reg  ( .D(\ctrl/counter/w7 ), .SI(
        n1037), .SE(test_se), .CK(clock), .RN(n758), .Q(n762), .QN(n702) );
  TBUF_X2 product_in_tri2_64_ ( .A(1'b0), .EN(n1042), .Z(product_in[64]) );
  TBUF_X2 product_in_tri3_0_ ( .A(1'b0), .EN(n1041), .Z(product_in[0]) );
  TBUF_X2 product_in_tri2_0_ ( .A(1'b0), .EN(n1042), .Z(product_in[0]) );
  TBUF_X2 product_in_tri2_2_ ( .A(data_operandB[1]), .EN(n1042), .Z(
        product_in[2]) );
  TBUF_X2 product_in_tri3_42_ ( .A(1'b0), .EN(n1067), .Z(product_in[42]) );
  TBUF_X2 product_in_tri2_42_ ( .A(1'b0), .EN(n1060), .Z(product_in[42]) );
  TBUF_X2 product_in_tri3_40_ ( .A(1'b0), .EN(n1067), .Z(product_in[40]) );
  TBUF_X2 product_in_tri2_40_ ( .A(1'b0), .EN(n1060), .Z(product_in[40]) );
  TBUF_X2 product_in_tri3_36_ ( .A(1'b0), .EN(n1063), .Z(product_in[36]) );
  TBUF_X2 product_in_tri3_38_ ( .A(1'b0), .EN(n1063), .Z(product_in[38]) );
  TBUF_X2 product_in_tri2_36_ ( .A(1'b0), .EN(n1064), .Z(product_in[36]) );
  TBUF_X2 product_in_tri2_38_ ( .A(1'b0), .EN(n1064), .Z(product_in[38]) );
  TBUF_X2 product_in_tri2_63_ ( .A(1'b0), .EN(n1045), .Z(product_in[63]) );
  TBUF_X2 product_in_tri3_63_ ( .A(1'b0), .EN(n1067), .Z(product_in[63]) );
  TBUF_X2 product_in_tri3_48_ ( .A(1'b0), .EN(n1067), .Z(product_in[48]) );
  TBUF_X2 product_in_tri3_50_ ( .A(1'b0), .EN(n1067), .Z(product_in[50]) );
  TBUF_X2 product_in_tri3_56_ ( .A(1'b0), .EN(n1067), .Z(product_in[56]) );
  TBUF_X2 product_in_tri3_58_ ( .A(1'b0), .EN(n1063), .Z(product_in[58]) );
  TBUF_X2 product_in_tri2_48_ ( .A(1'b0), .EN(n1060), .Z(product_in[48]) );
  TBUF_X2 product_in_tri2_50_ ( .A(1'b0), .EN(n1060), .Z(product_in[50]) );
  TBUF_X2 product_in_tri2_56_ ( .A(1'b0), .EN(n1064), .Z(product_in[56]) );
  TBUF_X2 product_in_tri2_58_ ( .A(1'b0), .EN(n1064), .Z(product_in[58]) );
  TBUF_X2 product_in_tri3_44_ ( .A(1'b0), .EN(n1063), .Z(product_in[44]) );
  TBUF_X2 product_in_tri3_46_ ( .A(1'b0), .EN(n1063), .Z(product_in[46]) );
  TBUF_X2 product_in_tri3_52_ ( .A(1'b0), .EN(n1063), .Z(product_in[52]) );
  TBUF_X2 product_in_tri3_54_ ( .A(1'b0), .EN(n1063), .Z(product_in[54]) );
  TBUF_X2 product_in_tri2_44_ ( .A(1'b0), .EN(n1064), .Z(product_in[44]) );
  TBUF_X2 product_in_tri2_46_ ( .A(1'b0), .EN(n1064), .Z(product_in[46]) );
  TBUF_X2 product_in_tri2_52_ ( .A(1'b0), .EN(n1042), .Z(product_in[52]) );
  TBUF_X2 product_in_tri2_54_ ( .A(1'b0), .EN(n1042), .Z(product_in[54]) );
  TBUF_X2 product_in_tri3_34_ ( .A(1'b0), .EN(n1041), .Z(product_in[34]) );
  TBUF_X2 product_in_tri2_34_ ( .A(1'b0), .EN(n1042), .Z(product_in[34]) );
  TBUF_X2 product_in_tri2_32_ ( .A(data_operandB[31]), .EN(n1042), .Z(
        product_in[32]) );
  TBUF_X2 product_in_tri2_25_ ( .A(data_operandB[24]), .EN(n1060), .Z(
        product_in[25]) );
  TBUF_X2 product_in_tri2_7_ ( .A(data_operandB[6]), .EN(n1045), .Z(
        product_in[7]) );
  TBUF_X2 product_in_tri2_4_ ( .A(data_operandB[3]), .EN(n1045), .Z(
        product_in[4]) );
  TBUF_X2 product_in_tri2_12_ ( .A(data_operandB[11]), .EN(n1045), .Z(
        product_in[12]) );
  TBUF_X2 product_in_tri2_15_ ( .A(data_operandB[14]), .EN(n1045), .Z(
        product_in[15]) );
  TBUF_X2 product_in_tri2_16_ ( .A(data_operandB[15]), .EN(n1045), .Z(
        product_in[16]) );
  TBUF_X2 product_in_tri2_20_ ( .A(data_operandB[19]), .EN(n1052), .Z(
        product_in[20]) );
  TBUF_X2 product_in_tri2_8_ ( .A(data_operandB[7]), .EN(n1045), .Z(
        product_in[8]) );
  TBUF_X2 product_in_tri2_9_ ( .A(data_operandB[8]), .EN(n1045), .Z(
        product_in[9]) );
  TBUF_X2 product_in_tri2_10_ ( .A(data_operandB[9]), .EN(n1045), .Z(
        product_in[10]) );
  TBUF_X2 product_in_tri2_11_ ( .A(data_operandB[10]), .EN(n1045), .Z(
        product_in[11]) );
  TBUF_X2 product_in_tri2_14_ ( .A(data_operandB[13]), .EN(n1045), .Z(
        product_in[14]) );
  TBUF_X2 product_in_tri2_30_ ( .A(data_operandB[29]), .EN(n1052), .Z(
        product_in[30]) );
  TBUF_X2 product_in_tri2_5_ ( .A(data_operandB[4]), .EN(n1052), .Z(
        product_in[5]) );
  TBUF_X2 product_in_tri2_29_ ( .A(data_operandB[28]), .EN(n1052), .Z(
        product_in[29]) );
  TBUF_X2 product_in_tri2_28_ ( .A(data_operandB[27]), .EN(n1052), .Z(
        product_in[28]) );
  TBUF_X2 product_in_tri2_18_ ( .A(data_operandB[17]), .EN(n1052), .Z(
        product_in[18]) );
  TBUF_X2 product_in_tri2_19_ ( .A(data_operandB[18]), .EN(n1052), .Z(
        product_in[19]) );
  TBUF_X2 product_in_tri2_24_ ( .A(data_operandB[23]), .EN(n1052), .Z(
        product_in[24]) );
  TBUF_X2 product_in_tri2_27_ ( .A(data_operandB[26]), .EN(n1052), .Z(
        product_in[27]) );
  TBUF_X2 product_in_tri2_26_ ( .A(data_operandB[25]), .EN(n1060), .Z(
        product_in[26]) );
  TBUF_X2 product_in_tri2_13_ ( .A(data_operandB[12]), .EN(n1045), .Z(
        product_in[13]) );
  TBUF_X2 product_in_tri2_3_ ( .A(data_operandB[2]), .EN(n1042), .Z(
        product_in[3]) );
  TBUF_X2 product_in_tri2_6_ ( .A(data_operandB[5]), .EN(n1052), .Z(
        product_in[6]) );
  TBUF_X2 product_in_tri2_23_ ( .A(data_operandB[22]), .EN(n1052), .Z(
        product_in[23]) );
  TBUF_X2 product_in_tri2_22_ ( .A(data_operandB[21]), .EN(n1060), .Z(
        product_in[22]) );
  TBUF_X2 product_in_tri2_17_ ( .A(data_operandB[16]), .EN(n1052), .Z(
        product_in[17]) );
  TBUF_X2 product_in_tri2_21_ ( .A(data_operandB[20]), .EN(n1052), .Z(
        product_in[21]) );
  TBUF_X2 product_in_tri2_1_ ( .A(data_operandB[0]), .EN(n1045), .Z(
        product_in[1]) );
  TBUF_X2 product_in_tri3_39_ ( .A(1'b0), .EN(n1067), .Z(product_in[39]) );
  TBUF_X2 product_in_tri2_39_ ( .A(1'b0), .EN(n1060), .Z(product_in[39]) );
  TBUF_X2 product_in_tri3_37_ ( .A(1'b0), .EN(n1067), .Z(product_in[37]) );
  TBUF_X2 product_in_tri3_45_ ( .A(1'b0), .EN(n1067), .Z(product_in[45]) );
  TBUF_X2 product_in_tri3_47_ ( .A(1'b0), .EN(n1067), .Z(product_in[47]) );
  TBUF_X2 product_in_tri3_53_ ( .A(1'b0), .EN(n1067), .Z(product_in[53]) );
  TBUF_X2 product_in_tri2_37_ ( .A(1'b0), .EN(n1060), .Z(product_in[37]) );
  TBUF_X2 product_in_tri2_45_ ( .A(1'b0), .EN(n1060), .Z(product_in[45]) );
  TBUF_X2 product_in_tri2_47_ ( .A(1'b0), .EN(n1060), .Z(product_in[47]) );
  TBUF_X2 product_in_tri2_53_ ( .A(1'b0), .EN(n1060), .Z(product_in[53]) );
  TBUF_X2 product_in_tri3_41_ ( .A(1'b0), .EN(n1063), .Z(product_in[41]) );
  TBUF_X2 product_in_tri3_43_ ( .A(1'b0), .EN(n1063), .Z(product_in[43]) );
  TBUF_X2 product_in_tri3_49_ ( .A(1'b0), .EN(n1063), .Z(product_in[49]) );
  TBUF_X2 product_in_tri3_51_ ( .A(1'b0), .EN(n1063), .Z(product_in[51]) );
  TBUF_X2 product_in_tri2_41_ ( .A(1'b0), .EN(n1064), .Z(product_in[41]) );
  TBUF_X2 product_in_tri3_35_ ( .A(1'b0), .EN(n1063), .Z(product_in[35]) );
  TBUF_X2 product_in_tri2_35_ ( .A(1'b0), .EN(n1064), .Z(product_in[35]) );
  TBUF_X2 product_in_tri2_43_ ( .A(1'b0), .EN(n1064), .Z(product_in[43]) );
  TBUF_X2 product_in_tri2_49_ ( .A(1'b0), .EN(n1064), .Z(product_in[49]) );
  TBUF_X2 product_in_tri2_51_ ( .A(1'b0), .EN(n1064), .Z(product_in[51]) );
  TBUF_X2 product_in_tri3_33_ ( .A(1'b0), .EN(n1041), .Z(product_in[33]) );
  TBUF_X2 product_in_tri2_33_ ( .A(1'b0), .EN(n1042), .Z(product_in[33]) );
  TBUF_X2 product_in_tri2_31_ ( .A(data_operandB[30]), .EN(n1042), .Z(
        product_in[31]) );
  TBUF_X2 product_in_tri3_61_ ( .A(1'b0), .EN(n1067), .Z(product_in[61]) );
  TBUF_X2 product_in_tri2_61_ ( .A(1'b0), .EN(n1060), .Z(product_in[61]) );
  TBUF_X2 product_in_tri3_59_ ( .A(1'b0), .EN(n1041), .Z(product_in[59]) );
  TBUF_X2 product_in_tri2_59_ ( .A(1'b0), .EN(n1042), .Z(product_in[59]) );
  TBUF_X2 product_in_tri3_62_ ( .A(1'b0), .EN(n1041), .Z(product_in[62]) );
  TBUF_X2 product_in_tri2_62_ ( .A(1'b0), .EN(n1042), .Z(product_in[62]) );
  TBUF_X2 product_in_tri3_60_ ( .A(1'b0), .EN(n1063), .Z(product_in[60]) );
  TBUF_X2 product_in_tri2_60_ ( .A(1'b0), .EN(n1064), .Z(product_in[60]) );
  TBUF_X2 product_in_tri3_55_ ( .A(1'b0), .EN(n1067), .Z(product_in[55]) );
  TBUF_X2 product_in_tri2_55_ ( .A(1'b0), .EN(n1064), .Z(product_in[55]) );
  TBUF_X2 product_in_tri3_57_ ( .A(1'b0), .EN(n1041), .Z(product_in[57]) );
  TBUF_X2 product_in_tri2_57_ ( .A(1'b0), .EN(n1042), .Z(product_in[57]) );
  TBUF_X2 product_in_tri_0_ ( .A(product_out[2]), .EN(n1043), .Z(product_in[0]) );
  TBUF_X2 product_in_tri4_0_ ( .A(1'b0), .EN(n1044), .Z(product_in[0]) );
  TBUF_X2 product_in_tri4_2_ ( .A(n120), .EN(n1048), .Z(product_in[2]) );
  TBUF_X2 product_in_tri3_2_ ( .A(n745), .EN(n1049), .Z(product_in[2]) );
  TBUF_X2 product_in_tri_2_ ( .A(product_out[4]), .EN(n1050), .Z(product_in[2]) );
  TBUF_X2 product_in_tri4_32_ ( .A(product_out[31]), .EN(n1061), .Z(
        product_in[32]) );
  TBUF_X2 product_in_tri4_25_ ( .A(product_out[24]), .EN(n1061), .Z(
        product_in[25]) );
  TBUF_X2 product_in_tri_25_ ( .A(product_out[27]), .EN(n1059), .Z(
        product_in[25]) );
  TBUF_X2 product_in_tri4_7_ ( .A(product_out[6]), .EN(n1048), .Z(
        product_in[7]) );
  TBUF_X2 product_in_tri4_3_ ( .A(product_out[2]), .EN(n1048), .Z(
        product_in[3]) );
  TBUF_X2 product_in_tri4_8_ ( .A(product_out[7]), .EN(n1048), .Z(
        product_in[8]) );
  TBUF_X2 product_in_tri4_4_ ( .A(product_out[3]), .EN(n1048), .Z(
        product_in[4]) );
  TBUF_X2 product_in_tri4_9_ ( .A(product_out[8]), .EN(n1048), .Z(
        product_in[9]) );
  TBUF_X2 product_in_tri4_11_ ( .A(product_out[10]), .EN(n1048), .Z(
        product_in[11]) );
  TBUF_X2 product_in_tri4_12_ ( .A(product_out[11]), .EN(n1048), .Z(
        product_in[12]) );
  TBUF_X2 product_in_tri4_15_ ( .A(product_out[14]), .EN(n1053), .Z(
        product_in[15]) );
  TBUF_X2 product_in_tri4_16_ ( .A(product_out[15]), .EN(n1053), .Z(
        product_in[16]) );
  TBUF_X2 product_in_tri4_20_ ( .A(product_out[19]), .EN(n1053), .Z(
        product_in[20]) );
  TBUF_X2 product_in_tri4_10_ ( .A(product_out[9]), .EN(n1048), .Z(
        product_in[10]) );
  TBUF_X2 product_in_tri4_14_ ( .A(product_out[13]), .EN(n1053), .Z(
        product_in[14]) );
  TBUF_X2 product_in_tri4_30_ ( .A(product_out[29]), .EN(n1053), .Z(
        product_in[30]) );
  TBUF_X2 product_in_tri4_5_ ( .A(product_out[4]), .EN(n1053), .Z(
        product_in[5]) );
  TBUF_X2 product_in_tri4_29_ ( .A(product_out[28]), .EN(n1061), .Z(
        product_in[29]) );
  TBUF_X2 product_in_tri4_28_ ( .A(product_out[27]), .EN(n1061), .Z(
        product_in[28]) );
  TBUF_X2 product_in_tri4_24_ ( .A(product_out[23]), .EN(n1061), .Z(
        product_in[24]) );
  TBUF_X2 product_in_tri4_27_ ( .A(product_out[26]), .EN(n1061), .Z(
        product_in[27]) );
  TBUF_X2 product_in_tri4_26_ ( .A(product_out[25]), .EN(n1061), .Z(
        product_in[26]) );
  TBUF_X2 product_in_tri3_7_ ( .A(n213), .EN(n1041), .Z(product_in[7]) );
  TBUF_X2 product_in_tri_7_ ( .A(product_out[9]), .EN(n1056), .Z(product_in[7]) );
  TBUF_X2 product_in_tri3_8_ ( .A(n212), .EN(n1041), .Z(product_in[8]) );
  TBUF_X2 product_in_tri_8_ ( .A(product_out[10]), .EN(n1051), .Z(
        product_in[8]) );
  TBUF_X2 product_in_tri3_4_ ( .A(n743), .EN(n1041), .Z(product_in[4]) );
  TBUF_X2 product_in_tri_4_ ( .A(product_out[6]), .EN(n1051), .Z(product_in[4]) );
  TBUF_X2 product_in_tri_9_ ( .A(product_out[11]), .EN(n1046), .Z(
        product_in[9]) );
  TBUF_X2 product_in_tri_11_ ( .A(product_out[13]), .EN(n1046), .Z(
        product_in[11]) );
  TBUF_X2 product_in_tri_12_ ( .A(product_out[14]), .EN(n1046), .Z(
        product_in[12]) );
  TBUF_X2 product_in_tri_15_ ( .A(product_out[17]), .EN(n1046), .Z(
        product_in[15]) );
  TBUF_X2 product_in_tri_16_ ( .A(product_out[18]), .EN(n1046), .Z(
        product_in[16]) );
  TBUF_X2 product_in_tri_20_ ( .A(product_out[22]), .EN(n1046), .Z(
        product_in[20]) );
  TBUF_X2 product_in_tri4_18_ ( .A(product_out[17]), .EN(n1053), .Z(
        product_in[18]) );
  TBUF_X2 product_in_tri4_19_ ( .A(product_out[18]), .EN(n1053), .Z(
        product_in[19]) );
  TBUF_X2 product_in_tri4_22_ ( .A(product_out[21]), .EN(n1061), .Z(
        product_in[22]) );
  TBUF_X2 product_in_tri_10_ ( .A(product_out[12]), .EN(n1046), .Z(
        product_in[10]) );
  TBUF_X2 product_in_tri_14_ ( .A(product_out[16]), .EN(n1046), .Z(
        product_in[14]) );
  TBUF_X2 product_in_tri_30_ ( .A(product_out[32]), .EN(n1059), .Z(
        product_in[30]) );
  TBUF_X2 product_in_tri3_9_ ( .A(n210), .EN(n1057), .Z(product_in[9]) );
  TBUF_X2 product_in_tri3_5_ ( .A(n741), .EN(n1054), .Z(product_in[5]) );
  TBUF_X2 product_in_tri_5_ ( .A(product_out[7]), .EN(n1055), .Z(product_in[5]) );
  TBUF_X2 product_in_tri_29_ ( .A(product_out[31]), .EN(n1059), .Z(
        product_in[29]) );
  TBUF_X2 product_in_tri_28_ ( .A(product_out[30]), .EN(n1059), .Z(
        product_in[28]) );
  TBUF_X2 product_in_tri_24_ ( .A(product_out[26]), .EN(n1059), .Z(
        product_in[24]) );
  TBUF_X2 product_in_tri_27_ ( .A(product_out[29]), .EN(n1059), .Z(
        product_in[27]) );
  TBUF_X2 product_in_tri_26_ ( .A(product_out[28]), .EN(n1059), .Z(
        product_in[26]) );
  TBUF_X2 product_in_tri4_6_ ( .A(product_out[5]), .EN(n1053), .Z(
        product_in[6]) );
  TBUF_X2 product_in_tri4_23_ ( .A(product_out[22]), .EN(n1061), .Z(
        product_in[23]) );
  TBUF_X2 product_in_tri_18_ ( .A(product_out[20]), .EN(n1046), .Z(
        product_in[18]) );
  TBUF_X2 product_in_tri_19_ ( .A(product_out[21]), .EN(n1046), .Z(
        product_in[19]) );
  TBUF_X2 product_in_tri3_3_ ( .A(n739), .EN(n1049), .Z(product_in[3]) );
  TBUF_X2 product_in_tri4_13_ ( .A(product_out[12]), .EN(n1053), .Z(
        product_in[13]) );
  TBUF_X2 product_in_tri_13_ ( .A(product_out[15]), .EN(n1046), .Z(
        product_in[13]) );
  TBUF_X2 product_in_tri3_6_ ( .A(n214), .EN(n1054), .Z(product_in[6]) );
  TBUF_X2 product_in_tri_6_ ( .A(product_out[8]), .EN(n1055), .Z(product_in[6]) );
  TBUF_X2 product_in_tri_23_ ( .A(product_out[25]), .EN(n1059), .Z(
        product_in[23]) );
  TBUF_X2 product_in_tri_22_ ( .A(product_out[24]), .EN(n1059), .Z(
        product_in[22]) );
  TBUF_X2 product_in_tri_3_ ( .A(product_out[5]), .EN(n1050), .Z(product_in[3]) );
  TBUF_X2 product_in_tri4_17_ ( .A(product_out[16]), .EN(n1053), .Z(
        product_in[17]) );
  TBUF_X2 product_in_tri4_21_ ( .A(product_out[20]), .EN(n1053), .Z(
        product_in[21]) );
  TBUF_X2 product_in_tri_17_ ( .A(product_out[19]), .EN(n1046), .Z(
        product_in[17]) );
  TBUF_X2 product_in_tri_21_ ( .A(product_out[23]), .EN(n1059), .Z(
        product_in[21]) );
  TBUF_X2 product_in_tri3_1_ ( .A(n747), .EN(n1041), .Z(product_in[1]) );
  TBUF_X2 product_in_tri_1_ ( .A(product_out[3]), .EN(n1046), .Z(product_in[1]) );
  TBUF_X2 product_in_tri4_31_ ( .A(product_out[30]), .EN(n1061), .Z(
        product_in[31]) );
  TBUF_X2 product_in_tri4_42_ ( .A(adder_out[9]), .EN(n1065), .Z(
        product_in[42]) );
  TBUF_X2 product_in_tri_42_ ( .A(adder_out[11]), .EN(n1066), .Z(
        product_in[42]) );
  TBUF_X2 product_in_tri_40_ ( .A(adder_out[9]), .EN(n1059), .Z(product_in[40]) );
  TBUF_X2 product_in_tri4_40_ ( .A(adder_out[7]), .EN(n1069), .Z(
        product_in[40]) );
  TBUF_X2 product_in_tri4_36_ ( .A(adder_out[3]), .EN(n1065), .Z(
        product_in[36]) );
  TBUF_X2 product_in_tri4_38_ ( .A(adder_out[5]), .EN(n1068), .Z(
        product_in[38]) );
  TBUF_X2 product_in_tri_36_ ( .A(adder_out[5]), .EN(n1066), .Z(product_in[36]) );
  TBUF_X2 product_in_tri_38_ ( .A(adder_out[7]), .EN(n1066), .Z(product_in[38]) );
  TBUF_X2 product_in_tri_34_ ( .A(adder_out[3]), .EN(n1043), .Z(product_in[34]) );
  TBUF_X2 product_in_tri4_44_ ( .A(adder_out[11]), .EN(n1068), .Z(
        product_in[44]) );
  TBUF_X2 product_in_tri4_46_ ( .A(adder_out[13]), .EN(n1068), .Z(
        product_in[46]) );
  TBUF_X2 product_in_tri_44_ ( .A(adder_out[13]), .EN(n1066), .Z(
        product_in[44]) );
  TBUF_X2 product_in_tri4_34_ ( .A(adder_out[1]), .EN(n1047), .Z(
        product_in[34]) );
  TBUF_X2 product_in_tri_32_ ( .A(adder_out[1]), .EN(n1043), .Z(product_in[32]) );
  TBUF_X2 product_in_tri3_32_ ( .A(n187), .EN(n1062), .Z(product_in[32]) );
  TBUF_X2 product_in_tri3_25_ ( .A(n708), .EN(n1062), .Z(product_in[25]) );
  TBUF_X2 product_in_tri3_16_ ( .A(n727), .EN(n1057), .Z(product_in[16]) );
  TBUF_X2 product_in_tri3_15_ ( .A(n729), .EN(n1058), .Z(product_in[15]) );
  TBUF_X2 product_in_tri3_11_ ( .A(n735), .EN(n1057), .Z(product_in[11]) );
  TBUF_X2 product_in_tri3_12_ ( .A(n733), .EN(n1057), .Z(product_in[12]) );
  TBUF_X2 product_in_tri3_20_ ( .A(n719), .EN(n1057), .Z(product_in[20]) );
  TBUF_X2 product_in_tri3_14_ ( .A(n731), .EN(n1058), .Z(product_in[14]) );
  TBUF_X2 product_in_tri3_10_ ( .A(n209), .EN(n1057), .Z(product_in[10]) );
  TBUF_X2 product_in_tri3_30_ ( .A(n704), .EN(n1062), .Z(product_in[30]) );
  TBUF_X2 product_in_tri3_29_ ( .A(n706), .EN(n1062), .Z(product_in[29]) );
  TBUF_X2 product_in_tri3_28_ ( .A(n713), .EN(n1062), .Z(product_in[28]) );
  TBUF_X2 product_in_tri3_24_ ( .A(n717), .EN(n1062), .Z(product_in[24]) );
  TBUF_X2 product_in_tri3_27_ ( .A(n710), .EN(n1062), .Z(product_in[27]) );
  TBUF_X2 product_in_tri3_26_ ( .A(n715), .EN(n1062), .Z(product_in[26]) );
  TBUF_X2 product_in_tri3_18_ ( .A(n723), .EN(n1057), .Z(product_in[18]) );
  TBUF_X2 product_in_tri3_19_ ( .A(n721), .EN(n1057), .Z(product_in[19]) );
  TBUF_X2 product_in_tri3_13_ ( .A(n737), .EN(n1058), .Z(product_in[13]) );
  TBUF_X2 product_in_tri3_23_ ( .A(n196), .EN(n1057), .Z(product_in[23]) );
  TBUF_X2 product_in_tri3_22_ ( .A(n197), .EN(n1062), .Z(product_in[22]) );
  TBUF_X2 product_in_tri3_17_ ( .A(n725), .EN(n1057), .Z(product_in[17]) );
  TBUF_X2 product_in_tri3_21_ ( .A(n198), .EN(n1057), .Z(product_in[21]) );
  TBUF_X2 product_in_tri4_33_ ( .A(adder_out[0]), .EN(n1048), .Z(
        product_in[33]) );
  TBUF_X2 product_in_tri_31_ ( .A(adder_out[0]), .EN(n1043), .Z(product_in[31]) );
  TBUF_X2 product_in_tri_33_ ( .A(adder_out[2]), .EN(n1056), .Z(product_in[33]) );
  TBUF_X2 product_in_tri_39_ ( .A(adder_out[8]), .EN(n1059), .Z(product_in[39]) );
  TBUF_X2 product_in_tri4_39_ ( .A(adder_out[6]), .EN(n1069), .Z(
        product_in[39]) );
  TBUF_X2 product_in_tri4_45_ ( .A(adder_out[12]), .EN(n1065), .Z(
        product_in[45]) );
  TBUF_X2 product_in_tri4_47_ ( .A(adder_out[14]), .EN(n1065), .Z(
        product_in[47]) );
  TBUF_X2 product_in_tri_45_ ( .A(adder_out[14]), .EN(n1066), .Z(
        product_in[45]) );
  TBUF_X2 product_in_tri4_41_ ( .A(adder_out[8]), .EN(n1065), .Z(
        product_in[41]) );
  TBUF_X2 product_in_tri4_43_ ( .A(adder_out[10]), .EN(n1065), .Z(
        product_in[43]) );
  TBUF_X2 product_in_tri_41_ ( .A(adder_out[10]), .EN(n1066), .Z(
        product_in[41]) );
  TBUF_X2 product_in_tri4_37_ ( .A(adder_out[4]), .EN(n1061), .Z(
        product_in[37]) );
  TBUF_X2 product_in_tri_37_ ( .A(adder_out[6]), .EN(n1066), .Z(product_in[37]) );
  TBUF_X2 product_in_tri4_35_ ( .A(adder_out[2]), .EN(n1065), .Z(
        product_in[35]) );
  TBUF_X2 product_in_tri_35_ ( .A(adder_out[4]), .EN(n1066), .Z(product_in[35]) );
  TBUF_X2 product_in_tri_43_ ( .A(adder_out[12]), .EN(n1066), .Z(
        product_in[43]) );
  TBUF_X2 product_in_tri3_31_ ( .A(n397), .EN(n1062), .Z(product_in[31]) );
  TBUF_X2 product_in_tri4_63_ ( .A(adder_out[30]), .EN(n1048), .Z(
        product_in[63]) );
  TBUF_X2 product_in_tri4_48_ ( .A(adder_out[15]), .EN(n1065), .Z(
        product_in[48]) );
  TBUF_X2 product_in_tri4_50_ ( .A(adder_out[17]), .EN(n1065), .Z(
        product_in[50]) );
  TBUF_X2 product_in_tri_48_ ( .A(adder_out[17]), .EN(n1066), .Z(
        product_in[48]) );
  TBUF_X2 product_in_tri_50_ ( .A(adder_out[19]), .EN(n1066), .Z(
        product_in[50]) );
  TBUF_X2 product_in_tri_46_ ( .A(adder_out[15]), .EN(n1066), .Z(
        product_in[46]) );
  TBUF_X2 product_in_tri4_52_ ( .A(adder_out[19]), .EN(n1068), .Z(
        product_in[52]) );
  TBUF_X2 product_in_tri4_56_ ( .A(adder_out[23]), .EN(n1068), .Z(
        product_in[56]) );
  TBUF_X2 product_in_tri4_58_ ( .A(adder_out[25]), .EN(n1068), .Z(
        product_in[58]) );
  TBUF_X2 product_in_tri_56_ ( .A(adder_out[25]), .EN(n1050), .Z(
        product_in[56]) );
  TBUF_X2 product_in_tri_58_ ( .A(adder_out[27]), .EN(n1050), .Z(
        product_in[58]) );
  TBUF_X2 product_in_tri4_54_ ( .A(adder_out[21]), .EN(n1070), .Z(
        product_in[54]) );
  TBUF_X2 product_in_tri_52_ ( .A(adder_out[21]), .EN(n1050), .Z(
        product_in[52]) );
  TBUF_X2 product_in_tri_54_ ( .A(adder_out[23]), .EN(n1050), .Z(
        product_in[54]) );
  TBUF_X2 product_in_tri4_1_ ( .A(n748), .EN(n1047), .Z(product_in[1]) );
  TBUF_X2 product_in_tri_47_ ( .A(adder_out[16]), .EN(n1066), .Z(
        product_in[47]) );
  TBUF_X2 product_in_tri4_53_ ( .A(adder_out[20]), .EN(n1065), .Z(
        product_in[53]) );
  TBUF_X2 product_in_tri4_49_ ( .A(adder_out[16]), .EN(n1068), .Z(
        product_in[49]) );
  TBUF_X2 product_in_tri4_51_ ( .A(adder_out[18]), .EN(n1068), .Z(
        product_in[51]) );
  TBUF_X2 product_in_tri_49_ ( .A(adder_out[18]), .EN(n1066), .Z(
        product_in[49]) );
  TBUF_X2 product_in_tri_51_ ( .A(adder_out[20]), .EN(n1066), .Z(
        product_in[51]) );
  TBUF_X2 product_in_tri_53_ ( .A(adder_out[22]), .EN(n1050), .Z(
        product_in[53]) );
  TBUF_X2 product_in_tri4_61_ ( .A(adder_out[28]), .EN(n1068), .Z(
        product_in[61]) );
  TBUF_X2 product_in_tri_61_ ( .A(adder_out[30]), .EN(n1050), .Z(
        product_in[61]) );
  TBUF_X2 product_in_tri4_59_ ( .A(adder_out[26]), .EN(n1070), .Z(
        product_in[59]) );
  TBUF_X2 product_in_tri_59_ ( .A(adder_out[28]), .EN(n1050), .Z(
        product_in[59]) );
  TBUF_X2 product_in_tri4_60_ ( .A(adder_out[27]), .EN(n1070), .Z(
        product_in[60]) );
  TBUF_X2 product_in_tri_60_ ( .A(adder_out[29]), .EN(n1050), .Z(
        product_in[60]) );
  TBUF_X2 product_in_tri4_55_ ( .A(adder_out[22]), .EN(n1068), .Z(
        product_in[55]) );
  TBUF_X2 product_in_tri_55_ ( .A(adder_out[24]), .EN(n1050), .Z(
        product_in[55]) );
  TBUF_X2 product_in_tri4_57_ ( .A(adder_out[24]), .EN(n1070), .Z(
        product_in[57]) );
  TBUF_X2 product_in_tri_57_ ( .A(adder_out[26]), .EN(n1050), .Z(
        product_in[57]) );
  TBUF_X2 product_in_tri_64_ ( .A(n625), .EN(n1050), .Z(product_in[64]) );
  TBUF_X2 product_in_tri_63_ ( .A(n625), .EN(n1056), .Z(product_in[63]) );
  TBUF_X2 product_in_tri_62_ ( .A(n71), .EN(n1059), .Z(product_in[62]) );
  TBUF_X2 product_in_tri4_62_ ( .A(adder_out[29]), .EN(n1071), .Z(
        product_in[62]) );
  SDFF_X1 \ctrl/cur_mult/q_reg  ( .D(\ctrl/cur_mult/n1 ), .SI(n117), .SE(
        test_se), .CK(clock), .Q(\ctrl/op_mult_int ), .QN(n116) );
  SDFF_X1 \ctrl/cur_div/q_reg  ( .D(\ctrl/cur_div/n1 ), .SI(n702), .SE(test_se), .CK(clock), .Q(\ctrl/op_div_int ), .QN(n117) );
  SDFF_X1 \product_reg/memory_32__dff/q_reg  ( .D(
        \product_reg/memory_32__dff/n1 ), .SI(product_out[31]), .SE(test_se), 
        .CK(clock), .Q(product_out[32]), .QN(n135) );
  SDFF_X1 \product_reg/memory_3__dff/q_reg  ( .D(
        \product_reg/memory_3__dff/n1 ), .SI(\product_reg/memory_2__dff/n7 ), 
        .SE(test_se), .CK(clock), .Q(product_out[3]), .QN(
        \product_reg/memory_3__dff/n5 ) );
  SDFF_X1 \product_reg/memory_4__dff/q_reg  ( .D(
        \product_reg/memory_4__dff/n1 ), .SI(product_out[3]), .SE(test_se), 
        .CK(clock), .Q(product_out[4]), .QN(\product_reg/memory_4__dff/n5 ) );
  SDFF_X1 \product_reg/memory_5__dff/q_reg  ( .D(
        \product_reg/memory_5__dff/n1 ), .SI(product_out[4]), .SE(test_se), 
        .CK(clock), .Q(product_out[5]), .QN(\product_reg/memory_5__dff/n5 ) );
  SDFF_X1 \product_reg/memory_6__dff/q_reg  ( .D(
        \product_reg/memory_6__dff/n1 ), .SI(product_out[5]), .SE(test_se), 
        .CK(clock), .Q(product_out[6]), .QN(\product_reg/memory_6__dff/n5 ) );
  SDFF_X1 \product_reg/memory_7__dff/q_reg  ( .D(
        \product_reg/memory_7__dff/n1 ), .SI(\product_reg/memory_6__dff/n5 ), 
        .SE(test_se), .CK(clock), .Q(product_out[7]), .QN(
        \product_reg/memory_7__dff/n5 ) );
  SDFF_X1 \product_reg/memory_8__dff/q_reg  ( .D(
        \product_reg/memory_8__dff/n1 ), .SI(product_out[7]), .SE(test_se), 
        .CK(clock), .Q(product_out[8]), .QN(\product_reg/memory_8__dff/n5 ) );
  SDFF_X1 \product_reg/memory_9__dff/q_reg  ( .D(
        \product_reg/memory_9__dff/n1 ), .SI(product_out[8]), .SE(test_se), 
        .CK(clock), .Q(product_out[9]), .QN(\product_reg/memory_9__dff/n5 ) );
  SDFF_X1 \product_reg/memory_10__dff/q_reg  ( .D(
        \product_reg/memory_10__dff/n1 ), .SI(\product_reg/memory_9__dff/n5 ), 
        .SE(test_se), .CK(clock), .Q(product_out[10]), .QN(
        \product_reg/memory_10__dff/n5 ) );
  SDFF_X1 \product_reg/memory_11__dff/q_reg  ( .D(
        \product_reg/memory_11__dff/n1 ), .SI(product_out[10]), .SE(test_se), 
        .CK(clock), .Q(product_out[11]), .QN(\product_reg/memory_11__dff/n5 )
         );
  SDFF_X1 \product_reg/memory_12__dff/q_reg  ( .D(
        \product_reg/memory_12__dff/n1 ), .SI(product_out[11]), .SE(test_se), 
        .CK(clock), .Q(product_out[12]), .QN(\product_reg/memory_12__dff/n5 )
         );
  SDFF_X1 \product_reg/memory_13__dff/q_reg  ( .D(
        \product_reg/memory_13__dff/n1 ), .SI(product_out[12]), .SE(test_se), 
        .CK(clock), .Q(product_out[13]), .QN(\product_reg/memory_13__dff/n5 )
         );
  SDFF_X1 \product_reg/memory_14__dff/q_reg  ( .D(
        \product_reg/memory_14__dff/n1 ), .SI(product_out[13]), .SE(test_se), 
        .CK(clock), .Q(product_out[14]), .QN(\product_reg/memory_14__dff/n5 )
         );
  SDFF_X1 \product_reg/memory_15__dff/q_reg  ( .D(
        \product_reg/memory_15__dff/n1 ), .SI(product_out[14]), .SE(test_se), 
        .CK(clock), .Q(product_out[15]), .QN(\product_reg/memory_15__dff/n5 )
         );
  SDFF_X1 \product_reg/memory_16__dff/q_reg  ( .D(
        \product_reg/memory_16__dff/n1 ), .SI(product_out[15]), .SE(test_se), 
        .CK(clock), .Q(product_out[16]), .QN(\product_reg/memory_16__dff/n5 )
         );
  SDFF_X1 \product_reg/memory_17__dff/q_reg  ( .D(
        \product_reg/memory_17__dff/n1 ), .SI(product_out[16]), .SE(test_se), 
        .CK(clock), .Q(product_out[17]), .QN(\product_reg/memory_17__dff/n5 )
         );
  SDFF_X1 \product_reg/memory_18__dff/q_reg  ( .D(
        \product_reg/memory_18__dff/n1 ), .SI(product_out[17]), .SE(test_se), 
        .CK(clock), .Q(product_out[18]), .QN(\product_reg/memory_18__dff/n5 )
         );
  SDFF_X1 \product_reg/memory_19__dff/q_reg  ( .D(
        \product_reg/memory_19__dff/n1 ), .SI(product_out[18]), .SE(test_se), 
        .CK(clock), .Q(product_out[19]), .QN(\product_reg/memory_19__dff/n5 )
         );
  SDFF_X1 \product_reg/memory_25__dff/q_reg  ( .D(
        \product_reg/memory_25__dff/n1 ), .SI(product_out[24]), .SE(test_se), 
        .CK(clock), .Q(product_out[25]), .QN(\product_reg/memory_25__dff/n5 )
         );
  SDFF_X1 \product_reg/memory_20__dff/q_reg  ( .D(
        \product_reg/memory_20__dff/n1 ), .SI(product_out[19]), .SE(test_se), 
        .CK(clock), .Q(product_out[20]), .QN(\product_reg/memory_20__dff/n5 )
         );
  SDFF_X1 \product_reg/memory_21__dff/q_reg  ( .D(
        \product_reg/memory_21__dff/n1 ), .SI(product_out[20]), .SE(test_se), 
        .CK(clock), .Q(product_out[21]), .QN(\product_reg/memory_21__dff/n5 )
         );
  SDFF_X1 \product_reg/memory_22__dff/q_reg  ( .D(
        \product_reg/memory_22__dff/n1 ), .SI(product_out[21]), .SE(test_se), 
        .CK(clock), .Q(product_out[22]), .QN(\product_reg/memory_22__dff/n5 )
         );
  SDFF_X1 \product_reg/memory_23__dff/q_reg  ( .D(
        \product_reg/memory_23__dff/n1 ), .SI(product_out[22]), .SE(test_se), 
        .CK(clock), .Q(product_out[23]), .QN(\product_reg/memory_23__dff/n5 )
         );
  SDFF_X1 \product_reg/memory_26__dff/q_reg  ( .D(
        \product_reg/memory_26__dff/n1 ), .SI(product_out[25]), .SE(test_se), 
        .CK(clock), .Q(product_out[26]), .QN(\product_reg/memory_26__dff/n5 )
         );
  SDFF_X1 \product_reg/memory_27__dff/q_reg  ( .D(
        \product_reg/memory_27__dff/n1 ), .SI(product_out[26]), .SE(test_se), 
        .CK(clock), .Q(product_out[27]), .QN(\product_reg/memory_27__dff/n5 )
         );
  SDFF_X1 \product_reg/memory_24__dff/q_reg  ( .D(
        \product_reg/memory_24__dff/n1 ), .SI(product_out[23]), .SE(test_se), 
        .CK(clock), .Q(product_out[24]), .QN(\product_reg/memory_24__dff/n5 )
         );
  SDFF_X1 \product_reg/memory_28__dff/q_reg  ( .D(
        \product_reg/memory_28__dff/n1 ), .SI(product_out[27]), .SE(test_se), 
        .CK(clock), .Q(product_out[28]), .QN(\product_reg/memory_28__dff/n5 )
         );
  SDFF_X1 \product_reg/memory_29__dff/q_reg  ( .D(
        \product_reg/memory_29__dff/n1 ), .SI(product_out[28]), .SE(test_se), 
        .CK(clock), .Q(product_out[29]), .QN(\product_reg/memory_29__dff/n5 )
         );
  SDFF_X1 \product_reg/memory_30__dff/q_reg  ( .D(
        \product_reg/memory_30__dff/n1 ), .SI(product_out[29]), .SE(test_se), 
        .CK(clock), .Q(product_out[30]), .QN(\product_reg/memory_30__dff/n5 )
         );
  SDFF_X1 \product_reg/memory_31__dff/q_reg  ( .D(
        \product_reg/memory_31__dff/n1 ), .SI(test_si3), .SE(test_se), .CK(
        clock), .Q(product_out[31]), .QN(\product_reg/memory_31__dff/n5 ) );
  SDFF_X1 \product_reg/memory_0__dff/q_reg  ( .D(n65), .SI(n116), .SE(test_se), 
        .CK(clock), .Q(n118), .QN(\product_reg/memory_0__dff/n5 ) );
  SDFF_X1 \product_reg/memory_33__dff/q_reg  ( .D(
        \product_reg/memory_33__dff/n1 ), .SI(product_out[32]), .SE(test_se), 
        .CK(clock), .Q(n1035), .QN(\product_reg/memory_33__dff/n5 ) );
  SDFF_X1 \product_reg/memory_34__dff/q_reg  ( .D(
        \product_reg/memory_34__dff/n1 ), .SI(n1035), .SE(test_se), .CK(clock), 
        .Q(n1034), .QN(\product_reg/memory_34__dff/n5 ) );
  SDFF_X1 \product_reg/memory_35__dff/q_reg  ( .D(
        \product_reg/memory_35__dff/n1 ), .SI(n1034), .SE(test_se), .CK(clock), 
        .Q(n1033), .QN(\product_reg/memory_35__dff/n5 ) );
  SDFF_X1 \product_reg/memory_36__dff/q_reg  ( .D(
        \product_reg/memory_36__dff/n1 ), .SI(n1033), .SE(test_se), .CK(clock), 
        .Q(n1032), .QN(\product_reg/memory_36__dff/n5 ) );
  SDFF_X1 \product_reg/memory_37__dff/q_reg  ( .D(
        \product_reg/memory_37__dff/n1 ), .SI(n1032), .SE(test_se), .CK(clock), 
        .Q(n1031), .QN(\product_reg/memory_37__dff/n5 ) );
  SDFF_X1 \product_reg/memory_38__dff/q_reg  ( .D(
        \product_reg/memory_38__dff/n1 ), .SI(n1031), .SE(test_se), .CK(clock), 
        .Q(n1030), .QN(\product_reg/memory_38__dff/n5 ) );
  SDFF_X1 \product_reg/memory_39__dff/q_reg  ( .D(
        \product_reg/memory_39__dff/n1 ), .SI(n1030), .SE(test_se), .CK(clock), 
        .Q(n1029), .QN(\product_reg/memory_39__dff/n5 ) );
  SDFF_X1 \product_reg/memory_40__dff/q_reg  ( .D(
        \product_reg/memory_40__dff/n1 ), .SI(n1029), .SE(test_se), .CK(clock), 
        .Q(n1028), .QN(\product_reg/memory_40__dff/n5 ) );
  SDFF_X1 \product_reg/memory_41__dff/q_reg  ( .D(
        \product_reg/memory_41__dff/n1 ), .SI(n1028), .SE(test_se), .CK(clock), 
        .Q(n1027), .QN(\product_reg/memory_41__dff/n5 ) );
  SDFF_X1 \product_reg/memory_42__dff/q_reg  ( .D(
        \product_reg/memory_42__dff/n1 ), .SI(n1027), .SE(test_se), .CK(clock), 
        .Q(n1026), .QN(\product_reg/memory_42__dff/n5 ) );
  SDFF_X1 \product_reg/memory_43__dff/q_reg  ( .D(
        \product_reg/memory_43__dff/n1 ), .SI(n1026), .SE(test_se), .CK(clock), 
        .Q(n1025), .QN(\product_reg/memory_43__dff/n5 ) );
  SDFF_X1 \product_reg/memory_44__dff/q_reg  ( .D(
        \product_reg/memory_44__dff/n1 ), .SI(n1025), .SE(test_se), .CK(clock), 
        .Q(n1024), .QN(\product_reg/memory_44__dff/n5 ) );
  SDFF_X1 \product_reg/memory_45__dff/q_reg  ( .D(
        \product_reg/memory_45__dff/n1 ), .SI(n1024), .SE(test_se), .CK(clock), 
        .Q(n1023), .QN(\product_reg/memory_45__dff/n5 ) );
  SDFF_X1 \product_reg/memory_46__dff/q_reg  ( .D(
        \product_reg/memory_46__dff/n1 ), .SI(n1023), .SE(test_se), .CK(clock), 
        .Q(n1022), .QN(\product_reg/memory_46__dff/n5 ) );
  SDFF_X1 \product_reg/memory_47__dff/q_reg  ( .D(
        \product_reg/memory_47__dff/n1 ), .SI(n1022), .SE(test_se), .CK(clock), 
        .Q(n1021), .QN(\product_reg/memory_47__dff/n5 ) );
  SDFF_X1 \product_reg/memory_48__dff/q_reg  ( .D(
        \product_reg/memory_48__dff/n1 ), .SI(n1021), .SE(test_se), .CK(clock), 
        .Q(n1020), .QN(\product_reg/memory_48__dff/n5 ) );
  SDFF_X1 \product_reg/memory_49__dff/q_reg  ( .D(
        \product_reg/memory_49__dff/n1 ), .SI(n1020), .SE(test_se), .CK(clock), 
        .Q(n1019), .QN(\product_reg/memory_49__dff/n5 ) );
  SDFF_X1 \product_reg/memory_50__dff/q_reg  ( .D(
        \product_reg/memory_50__dff/n1 ), .SI(n1019), .SE(test_se), .CK(clock), 
        .Q(n1018), .QN(\product_reg/memory_50__dff/n5 ) );
  SDFF_X1 \product_reg/memory_51__dff/q_reg  ( .D(
        \product_reg/memory_51__dff/n1 ), .SI(n1018), .SE(test_se), .CK(clock), 
        .Q(n1017), .QN(\product_reg/memory_51__dff/n5 ) );
  SDFF_X1 \product_reg/memory_52__dff/q_reg  ( .D(
        \product_reg/memory_52__dff/n1 ), .SI(n1017), .SE(test_se), .CK(clock), 
        .Q(n1016), .QN(\product_reg/memory_52__dff/n5 ) );
  SDFF_X1 \product_reg/memory_53__dff/q_reg  ( .D(
        \product_reg/memory_53__dff/n1 ), .SI(n1016), .SE(test_se), .CK(clock), 
        .Q(n1015), .QN(\product_reg/memory_53__dff/n5 ) );
  SDFF_X1 \product_reg/memory_54__dff/q_reg  ( .D(
        \product_reg/memory_54__dff/n1 ), .SI(n1015), .SE(test_se), .CK(clock), 
        .Q(n136), .QN(\product_reg/memory_54__dff/n5 ) );
  SDFF_X1 \product_reg/memory_56__dff/q_reg  ( .D(
        \product_reg/memory_56__dff/n1 ), .SI(n137), .SE(test_se), .CK(clock), 
        .Q(n1014), .QN(\product_reg/memory_56__dff/n5 ) );
  SDFF_X1 \product_reg/memory_55__dff/q_reg  ( .D(
        \product_reg/memory_55__dff/n1 ), .SI(n136), .SE(test_se), .CK(clock), 
        .Q(n137), .QN(\product_reg/memory_55__dff/n5 ) );
  SDFF_X1 \product_reg/memory_57__dff/q_reg  ( .D(
        \product_reg/memory_57__dff/n1 ), .SI(n1014), .SE(test_se), .CK(clock), 
        .Q(n1013), .QN(\product_reg/memory_57__dff/n5 ) );
  SDFF_X1 \product_reg/memory_58__dff/q_reg  ( .D(
        \product_reg/memory_58__dff/n1 ), .SI(n1013), .SE(test_se), .CK(clock), 
        .Q(n1012), .QN(\product_reg/memory_58__dff/n5 ) );
  SDFF_X1 \product_reg/memory_61__dff/q_reg  ( .D(
        \product_reg/memory_61__dff/n1 ), .SI(n1010), .SE(test_se), .CK(clock), 
        .Q(n1009), .QN(\product_reg/memory_61__dff/n5 ) );
  SDFF_X1 \product_reg/memory_59__dff/q_reg  ( .D(
        \product_reg/memory_59__dff/n1 ), .SI(n1012), .SE(test_se), .CK(clock), 
        .Q(n1011), .QN(\product_reg/memory_59__dff/n5 ) );
  SDFF_X1 \product_reg/memory_60__dff/q_reg  ( .D(
        \product_reg/memory_60__dff/n1 ), .SI(n1011), .SE(test_se), .CK(clock), 
        .Q(n1010), .QN(\product_reg/memory_60__dff/n5 ) );
  SDFF_X1 \product_reg/memory_62__dff/q_reg  ( .D(
        \product_reg/memory_62__dff/n1 ), .SI(n1009), .SE(test_se), .CK(clock), 
        .Q(n1008), .QN(\product_reg/memory_62__dff/n5 ) );
  SDFF_X1 \product_reg/memory_1__dff/q_reg  ( .D(
        \product_reg/memory_1__dff/n1 ), .SI(n118), .SE(test_se), .CK(clock), 
        .Q(n120), .QN(\product_reg/memory_1__dff/n8 ) );
  SDFF_X1 \product_reg/memory_64__dff/q_reg  ( .D(
        \product_reg/memory_64__dff/n1 ), .SI(n1007), .SE(test_se), .CK(clock), 
        .Q(test_so3), .QN(\product_reg/memory_64__dff/n5 ) );
  SDFF_X1 \product_reg/memory_63__dff/q_reg  ( .D(
        \product_reg/memory_63__dff/n1 ), .SI(n1008), .SE(test_se), .CK(clock), 
        .Q(n1007), .QN(\product_reg/memory_63__dff/n6 ) );
  SDFF_X1 \product_reg/memory_2__dff/q_reg  ( .D(n899), .SI(n120), .SE(test_se), .CK(clock), .Q(product_out[2]), .QN(\product_reg/memory_2__dff/n7 ) );
  NAND2_X2 U795 ( .A1(\ctrl/op_mult_int ), .A2(n758), .ZN(n760) );
  AND2_X4 U796 ( .A1(\ctrl/op_div_int ), .A2(n758), .ZN(n761) );
  INV_X4 U864 ( .A(n849), .ZN(n841) );
  INV_X4 U865 ( .A(n848), .ZN(n845) );
  INV_X4 U866 ( .A(n848), .ZN(n846) );
  INV_X4 U867 ( .A(n848), .ZN(n847) );
  INV_X4 U868 ( .A(n848), .ZN(n842) );
  INV_X4 U869 ( .A(n848), .ZN(n844) );
  INV_X4 U870 ( .A(n848), .ZN(n843) );
  INV_X4 U871 ( .A(n882), .ZN(n873) );
  INV_X4 U872 ( .A(n882), .ZN(n876) );
  INV_X4 U873 ( .A(n882), .ZN(n874) );
  INV_X4 U874 ( .A(n882), .ZN(n875) );
  INV_X4 U875 ( .A(n882), .ZN(n877) );
  INV_X4 U876 ( .A(n882), .ZN(n878) );
  INV_X4 U877 ( .A(n872), .ZN(n869) );
  INV_X4 U878 ( .A(n872), .ZN(n870) );
  OAI21_X2 U879 ( .B1(n672), .B2(n115), .A(n673), .ZN(n577) );
  AOI21_X2 U880 ( .B1(n87), .B2(n444), .A(n448), .ZN(n441) );
  AOI21_X2 U881 ( .B1(n510), .B2(n74), .A(n511), .ZN(n504) );
  OAI21_X2 U882 ( .B1(n427), .B2(n425), .A(n428), .ZN(n650) );
  AOI21_X2 U883 ( .B1(n555), .B2(n100), .A(n556), .ZN(n548) );
  AOI21_X2 U884 ( .B1(n624), .B2(n92), .A(n626), .ZN(n617) );
  AOI21_X2 U885 ( .B1(n85), .B2(n78), .A(n435), .ZN(n425) );
  AOI21_X2 U886 ( .B1(n97), .B2(n76), .A(n583), .ZN(n572) );
  AOI21_X2 U887 ( .B1(n89), .B2(n650), .A(n651), .ZN(n642) );
  AOI21_X2 U888 ( .B1(n96), .B2(n592), .A(n593), .ZN(n585) );
  AOI21_X2 U889 ( .B1(n523), .B2(n104), .A(n524), .ZN(n516) );
  OAI21_X2 U890 ( .B1(n600), .B2(n601), .A(n602), .ZN(n592) );
  OAI21_X2 U891 ( .B1(n563), .B2(n75), .A(n564), .ZN(n555) );
  OAI21_X2 U892 ( .B1(n633), .B2(n77), .A(n634), .ZN(n624) );
  OAI21_X2 U893 ( .B1(n504), .B2(n505), .A(n506), .ZN(n503) );
  OAI21_X2 U894 ( .B1(n443), .B2(n441), .A(n442), .ZN(n438) );
  OAI21_X2 U895 ( .B1(n490), .B2(n485), .A(n491), .ZN(n460) );
  OAI21_X2 U896 ( .B1(n572), .B2(n573), .A(n574), .ZN(n566) );
  OAI21_X2 U897 ( .B1(n642), .B2(n643), .A(n644), .ZN(n636) );
  OAI21_X2 U898 ( .B1(n547), .B2(n548), .A(n549), .ZN(n540) );
  OAI21_X2 U899 ( .B1(n616), .B2(n617), .A(n618), .ZN(n611) );
  INV_X4 U900 ( .A(n830), .ZN(n857) );
  INV_X4 U901 ( .A(n830), .ZN(n858) );
  INV_X4 U902 ( .A(n831), .ZN(n860) );
  INV_X4 U903 ( .A(n833), .ZN(n851) );
  INV_X4 U904 ( .A(n832), .ZN(n856) );
  NOR2_X2 U905 ( .A1(n557), .A2(n556), .ZN(n558) );
  NOR2_X2 U906 ( .A1(n465), .A2(n464), .ZN(n476) );
  NOR2_X2 U907 ( .A1(n594), .A2(n593), .ZN(n595) );
  NOR2_X2 U908 ( .A1(n525), .A2(n524), .ZN(n526) );
  NOR2_X2 U909 ( .A1(n547), .A2(n101), .ZN(n550) );
  NOR2_X2 U910 ( .A1(n573), .A2(n98), .ZN(n578) );
  INV_X4 U911 ( .A(n760), .ZN(n848) );
  INV_X4 U912 ( .A(n760), .ZN(n849) );
  INV_X4 U913 ( .A(n831), .ZN(n861) );
  INV_X4 U914 ( .A(n866), .ZN(n863) );
  INV_X4 U915 ( .A(n866), .ZN(n864) );
  INV_X4 U916 ( .A(n833), .ZN(n852) );
  INV_X4 U917 ( .A(n832), .ZN(n855) );
  INV_X4 U918 ( .A(n830), .ZN(n859) );
  INV_X4 U919 ( .A(n669), .ZN(n888) );
  INV_X4 U920 ( .A(n669), .ZN(n889) );
  INV_X4 U921 ( .A(n866), .ZN(n865) );
  NOR2_X2 U922 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X2 U923 ( .A1(n84), .A2(n427), .ZN(n426) );
  NOR2_X2 U924 ( .A1(n616), .A2(n93), .ZN(n619) );
  NOR2_X2 U925 ( .A1(n643), .A2(n90), .ZN(n645) );
  NOR2_X2 U926 ( .A1(n105), .A2(n112), .ZN(n511) );
  INV_X4 U927 ( .A(n831), .ZN(n862) );
  INV_X4 U928 ( .A(n832), .ZN(n854) );
  INV_X4 U929 ( .A(n833), .ZN(n853) );
  INV_X4 U930 ( .A(n669), .ZN(n887) );
  INV_X4 U931 ( .A(n216), .ZN(n880) );
  INV_X4 U932 ( .A(n216), .ZN(n879) );
  INV_X4 U933 ( .A(n216), .ZN(data_resultRDY) );
  INV_X4 U934 ( .A(n761), .ZN(n839) );
  INV_X4 U935 ( .A(n761), .ZN(n838) );
  INV_X4 U936 ( .A(n761), .ZN(n837) );
  INV_X4 U937 ( .A(n761), .ZN(n836) );
  INV_X4 U938 ( .A(n761), .ZN(n835) );
  INV_X4 U939 ( .A(n761), .ZN(n840) );
  INV_X4 U940 ( .A(n834), .ZN(n871) );
  INV_X4 U941 ( .A(ctrl_MULT), .ZN(n883) );
  INV_X4 U942 ( .A(ctrl_MULT), .ZN(n884) );
  INV_X4 U943 ( .A(ctrl_MULT), .ZN(n885) );
  INV_X4 U944 ( .A(ctrl_MULT), .ZN(n886) );
  INV_X4 U945 ( .A(n834), .ZN(n872) );
  NAND3_X2 U946 ( .A1(n108), .A2(n484), .A3(n72), .ZN(n493) );
  AOI21_X2 U947 ( .B1(n664), .B2(n451), .A(n456), .ZN(n444) );
  AOI21_X2 U948 ( .B1(n577), .B2(n666), .A(n667), .ZN(n485) );
  AOI21_X2 U949 ( .B1(n113), .B2(n82), .A(n576), .ZN(n667) );
  OAI21_X2 U950 ( .B1(n531), .B2(n532), .A(n533), .ZN(n523) );
  NOR2_X2 U951 ( .A1(n534), .A2(n535), .ZN(n531) );
  AOI21_X2 U952 ( .B1(n436), .B2(n439), .A(n79), .ZN(n429) );
  OAI21_X2 U953 ( .B1(n439), .B2(n436), .A(n438), .ZN(n661) );
  OAI21_X2 U954 ( .B1(n72), .B2(n481), .A(n482), .ZN(n463) );
  NOR2_X2 U955 ( .A1(n483), .A2(n484), .ZN(n481) );
  OAI21_X2 U956 ( .B1(n497), .B2(n73), .A(n498), .ZN(n496) );
  NOR2_X2 U957 ( .A1(n499), .A2(n500), .ZN(n497) );
  NOR2_X2 U958 ( .A1(n693), .A2(n694), .ZN(n672) );
  AND2_X2 U959 ( .A1(n691), .A2(n850), .ZN(n830) );
  AND2_X2 U960 ( .A1(n691), .A2(n847), .ZN(n831) );
  OR2_X2 U961 ( .A1(n691), .A2(n841), .ZN(n832) );
  OR2_X2 U962 ( .A1(n691), .A2(n848), .ZN(n833) );
  NOR2_X2 U963 ( .A1(n222), .A2(n841), .ZN(n625) );
  NOR2_X2 U964 ( .A1(n563), .A2(n99), .ZN(n565) );
  NOR2_X2 U965 ( .A1(n600), .A2(n95), .ZN(n603) );
  NOR2_X2 U966 ( .A1(n584), .A2(n583), .ZN(n586) );
  AOI21_X2 U967 ( .B1(n112), .B2(n105), .A(n511), .ZN(n517) );
  AOI21_X2 U968 ( .B1(n539), .B2(n538), .A(n541), .ZN(n544) );
  AOI21_X2 U969 ( .B1(n610), .B2(n609), .A(n612), .ZN(n613) );
  NAND3_X2 U970 ( .A1(n103), .A2(n535), .A3(n532), .ZN(n537) );
  NAND3_X2 U971 ( .A1(n107), .A2(n500), .A3(n73), .ZN(n502) );
  NOR2_X2 U972 ( .A1(n660), .A2(n659), .ZN(n427) );
  NOR2_X2 U973 ( .A1(n455), .A2(n454), .ZN(n456) );
  NOR2_X2 U974 ( .A1(n605), .A2(n606), .ZN(n600) );
  NOR2_X2 U975 ( .A1(n638), .A2(n639), .ZN(n633) );
  NOR2_X2 U976 ( .A1(n489), .A2(n488), .ZN(n490) );
  NOR2_X2 U977 ( .A1(n580), .A2(n579), .ZN(n573) );
  NOR2_X2 U978 ( .A1(n647), .A2(n646), .ZN(n643) );
  NOR2_X2 U979 ( .A1(n621), .A2(n620), .ZN(n616) );
  NOR2_X2 U980 ( .A1(n450), .A2(n449), .ZN(n447) );
  NOR2_X2 U981 ( .A1(n663), .A2(n662), .ZN(n443) );
  NOR2_X2 U982 ( .A1(n609), .A2(n610), .ZN(n612) );
  NOR2_X2 U983 ( .A1(n589), .A2(n588), .ZN(n584) );
  NOR2_X2 U984 ( .A1(n433), .A2(n432), .ZN(n434) );
  NOR2_X2 U985 ( .A1(n656), .A2(n655), .ZN(n652) );
  NOR2_X2 U986 ( .A1(n597), .A2(n596), .ZN(n594) );
  NOR2_X2 U987 ( .A1(n630), .A2(n629), .ZN(n627) );
  INV_X4 U988 ( .A(n868), .ZN(n866) );
  INV_X4 U989 ( .A(n760), .ZN(n850) );
  INV_X4 U990 ( .A(n868), .ZN(n867) );
  NOR3_X2 U991 ( .A1(n402), .A2(n401), .A3(n400), .ZN(n351) );
  NOR3_X2 U992 ( .A1(n408), .A2(n410), .A3(n411), .ZN(n413) );
  AOI21_X2 U993 ( .B1(n454), .B2(n455), .A(n456), .ZN(n452) );
  NOR2_X2 U994 ( .A1(n633), .A2(n91), .ZN(n635) );
  NOR2_X2 U995 ( .A1(n672), .A2(n83), .ZN(n690) );
  NOR2_X2 U996 ( .A1(n490), .A2(n88), .ZN(n486) );
  NOR2_X2 U997 ( .A1(n652), .A2(n651), .ZN(n653) );
  NOR2_X2 U998 ( .A1(n434), .A2(n435), .ZN(n430) );
  NOR3_X2 U999 ( .A1(n348), .A2(n302), .A3(n304), .ZN(n418) );
  NOR2_X2 U1000 ( .A1(n338), .A2(n339), .ZN(n407) );
  NOR2_X2 U1001 ( .A1(n319), .A2(n320), .ZN(n345) );
  NOR3_X2 U1002 ( .A1(n327), .A2(n328), .A3(n417), .ZN(n356) );
  NOR3_X2 U1003 ( .A1(n347), .A2(n348), .A3(n349), .ZN(n303) );
  NOR2_X2 U1004 ( .A1(n568), .A2(n569), .ZN(n563) );
  NOR2_X2 U1005 ( .A1(n552), .A2(n551), .ZN(n547) );
  NOR2_X2 U1006 ( .A1(n512), .A2(n513), .ZN(n505) );
  NOR2_X2 U1007 ( .A1(n538), .A2(n539), .ZN(n541) );
  NOR2_X2 U1008 ( .A1(n528), .A2(n527), .ZN(n525) );
  NOR2_X2 U1009 ( .A1(n560), .A2(n559), .ZN(n557) );
  NOR2_X2 U1010 ( .A1(n478), .A2(n477), .ZN(n465) );
  NAND3_X2 U1011 ( .A1(n129), .A2(n128), .A3(n413), .ZN(n400) );
  NAND3_X2 U1012 ( .A1(n124), .A2(n346), .A3(n345), .ZN(n342) );
  NOR2_X2 U1013 ( .A1(n356), .A2(n119), .ZN(n337) );
  OAI21_X2 U1014 ( .B1(n328), .B2(n327), .A(n417), .ZN(n416) );
  NOR2_X2 U1015 ( .A1(n316), .A2(n317), .ZN(n323) );
  NOR2_X2 U1016 ( .A1(n342), .A2(n343), .ZN(n341) );
  OAI21_X2 U1017 ( .B1(n444), .B2(n445), .A(n446), .ZN(adder_out[5]) );
  OAI21_X2 U1018 ( .B1(n447), .B2(n448), .A(n444), .ZN(n446) );
  NOR2_X2 U1019 ( .A1(n348), .A2(n349), .ZN(n350) );
  NAND3_X2 U1020 ( .A1(n130), .A2(n131), .A3(n351), .ZN(n349) );
  NOR2_X2 U1021 ( .A1(n401), .A2(n400), .ZN(n403) );
  NAND3_X2 U1022 ( .A1(n126), .A2(n127), .A3(n407), .ZN(n411) );
  NOR2_X2 U1023 ( .A1(n410), .A2(n411), .ZN(n409) );
  NOR2_X2 U1024 ( .A1(n337), .A2(n897), .ZN(n187) );
  OAI21_X2 U1025 ( .B1(n116), .B2(n424), .A(n886), .ZN(\ctrl/cur_mult/n1 ) );
  AND2_X2 U1026 ( .A1(n366), .A2(n762), .ZN(n834) );
  OAI21_X2 U1027 ( .B1(\product_reg/memory_1__dff/n8 ), .B2(
        \product_reg/memory_0__dff/n5 ), .A(product_out[2]), .ZN(n695) );
  AOI21_X2 U1028 ( .B1(n463), .B2(n109), .A(n464), .ZN(n462) );
  AOI21_X2 U1029 ( .B1(\product_reg/memory_1__dff/n8 ), .B2(n118), .A(
        ctrl_MULT), .ZN(n696) );
  INV_X4 U1030 ( .A(n468), .ZN(n868) );
  OAI21_X2 U1031 ( .B1(\product_reg/memory_0__dff/n5 ), .B2(n697), .A(n700), 
        .ZN(n699) );
  NAND3_X2 U1032 ( .A1(\product_reg/memory_1__dff/n8 ), .A2(product_out[2]), 
        .A3(\product_reg/memory_0__dff/n5 ), .ZN(n700) );
  INV_X4 U1033 ( .A(n216), .ZN(n882) );
  OAI21_X2 U1034 ( .B1(n117), .B2(n424), .A(n890), .ZN(\ctrl/cur_div/n1 ) );
  NOR2_X2 U1035 ( .A1(ctrl_DIV), .A2(ctrl_MULT), .ZN(n758) );
  AOI21_X2 U1036 ( .B1(n354), .B2(n355), .A(n356), .ZN(n353) );
  AOI222_X1 U1037 ( .A1(n138), .A2(data_result[31]), .B1(n365), .B2(n366), 
        .C1(n367), .C2(n368), .ZN(n352) );
  NAND3_X2 U1038 ( .A1(\product_reg/memory_63__dff/n6 ), .A2(n135), .A3(
        \product_reg/memory_62__dff/n5 ), .ZN(n388) );
  NOR2_X2 U1039 ( .A1(data_result[31]), .A2(n389), .ZN(n365) );
  INV_X4 U1040 ( .A(data_operandA[31]), .ZN(n897) );
  INV_X4 U1041 ( .A(ctrl_DIV), .ZN(n895) );
  INV_X4 U1042 ( .A(ctrl_DIV), .ZN(n896) );
  INV_X4 U1043 ( .A(data_operandA[31]), .ZN(n898) );
  INV_X4 U1044 ( .A(ctrl_DIV), .ZN(n890) );
  INV_X4 U1045 ( .A(ctrl_DIV), .ZN(n891) );
  INV_X4 U1046 ( .A(ctrl_DIV), .ZN(n893) );
  INV_X4 U1047 ( .A(ctrl_DIV), .ZN(n894) );
  INV_X4 U1048 ( .A(ctrl_DIV), .ZN(n892) );
  INV_X1 U1049 ( .A(n755), .ZN(n899) );
  NOR2_X1 U1133 ( .A1(test_se), .A2(n983), .ZN(n1050) );
  NAND2_X1 U1134 ( .A1(n984), .A2(n985), .ZN(n1042) );
  NOR2_X1 U1135 ( .A1(test_se), .A2(n986), .ZN(n1056) );
  NAND2_X1 U1136 ( .A1(n984), .A2(n987), .ZN(n1048) );
  NAND2_X1 U1137 ( .A1(n984), .A2(n988), .ZN(n1067) );
  NAND2_X1 U1138 ( .A1(n984), .A2(n989), .ZN(n1045) );
  NOR2_X1 U1139 ( .A1(test_se), .A2(n987), .ZN(n1071) );
  NAND2_X1 U1140 ( .A1(n984), .A2(n990), .ZN(n1059) );
  NAND2_X1 U1141 ( .A1(n984), .A2(n991), .ZN(n1041) );
  NAND2_X1 U1142 ( .A1(n984), .A2(n992), .ZN(n1068) );
  NAND2_X1 U1143 ( .A1(n984), .A2(n993), .ZN(n1060) );
  NAND2_X1 U1144 ( .A1(n984), .A2(n994), .ZN(n1070) );
  NAND2_X1 U1145 ( .A1(n984), .A2(n995), .ZN(n1064) );
  NAND2_X1 U1146 ( .A1(n984), .A2(n996), .ZN(n1063) );
  NAND2_X1 U1147 ( .A1(n984), .A2(n997), .ZN(n1065) );
  NOR2_X1 U1148 ( .A1(test_se), .A2(n998), .ZN(n1066) );
  NOR2_X1 U1149 ( .A1(test_se), .A2(n997), .ZN(n1069) );
  NAND2_X1 U1150 ( .A1(n984), .A2(n999), .ZN(n1061) );
  NOR2_X1 U1151 ( .A1(test_se), .A2(n992), .ZN(n1047) );
  NAND2_X1 U1152 ( .A1(n984), .A2(n986), .ZN(n1043) );
  NOR2_X1 U1153 ( .A1(test_se), .A2(n1000), .ZN(n1062) );
  NAND2_X1 U1154 ( .A1(n984), .A2(n1001), .ZN(n1053) );
  NAND2_X1 U1155 ( .A1(n984), .A2(n1002), .ZN(n1052) );
  NOR2_X1 U1156 ( .A1(test_se), .A2(n1003), .ZN(n1057) );
  NAND2_X1 U1157 ( .A1(n984), .A2(n1004), .ZN(n1046) );
  NOR2_X1 U1158 ( .A1(test_se), .A2(n991), .ZN(n1058) );
  NOR2_X1 U1159 ( .A1(test_se), .A2(n1004), .ZN(n1051) );
  NOR2_X1 U1160 ( .A1(test_se), .A2(n990), .ZN(n1055) );
  NAND2_X1 U1161 ( .A1(n984), .A2(n1003), .ZN(n1054) );
  NAND2_X1 U1162 ( .A1(n984), .A2(n1000), .ZN(n1049) );
  NOR2_X1 U1163 ( .A1(test_se), .A2(n999), .ZN(n1044) );
  INV_X1 U1164 ( .A(n837), .ZN(n999) );
  INV_X1 U1165 ( .A(n839), .ZN(n992) );
  INV_X1 U1166 ( .A(n841), .ZN(n983) );
  INV_X1 U1167 ( .A(n844), .ZN(n1004) );
  INV_X1 U1168 ( .A(n843), .ZN(n990) );
  INV_X1 U1169 ( .A(n845), .ZN(n986) );
  INV_X1 U1170 ( .A(n891), .ZN(n1003) );
  INV_X1 U1171 ( .A(n892), .ZN(n991) );
  INV_X1 U1172 ( .A(n890), .ZN(n1000) );
  INV_X1 U1173 ( .A(n842), .ZN(n998) );
  INV_X1 U1174 ( .A(n838), .ZN(n997) );
  INV_X1 U1175 ( .A(n835), .ZN(n987) );
  INV_X1 U1176 ( .A(test_se), .ZN(n984) );
  INV_X1 U1177 ( .A(n207), .ZN(n985) );
  INV_X1 U1178 ( .A(n894), .ZN(n988) );
  INV_X1 U1179 ( .A(n886), .ZN(n989) );
  INV_X1 U1180 ( .A(n884), .ZN(n993) );
  INV_X1 U1181 ( .A(n840), .ZN(n994) );
  INV_X1 U1182 ( .A(n883), .ZN(n995) );
  INV_X1 U1183 ( .A(n893), .ZN(n996) );
  INV_X1 U1184 ( .A(n836), .ZN(n1001) );
  INV_X1 U1185 ( .A(n885), .ZN(n1002) );
endmodule

