
module divider_dshift ( i_clk, i_rst, i_dividend, i_divisor, i_start, o_ready, 
        o_quotient, o_remainder );
  input [31:0] i_dividend;
  input [31:0] i_divisor;
  output [31:0] o_quotient;
  output [31:0] o_remainder;
  input i_clk, i_rst, i_start;
  output o_ready;
  wire   ready, reg_carry, n_1_net__3_, n_1_net__2_, n_1_net__1_, n_1_net__0_,
         state_reg_1_0, N264, N265, N266, N267, N268, N269, N270, N271, N272,
         N273, N274, N275, N276, N277, N278, N279, N280, N281, N282, N283,
         N284, N285, N286, N287, N288, N289, N290, N291, N292, N293, N294,
         N295, n701, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n829, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n870, n934, n935, n936, n937, n938, n939, n940, n941, n944,
         n945, n946, n947, n948, n949, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1113, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1296, n1297,
         n1350, n1769, n1770, n1771, n1772, n1773, n1829, n1864, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
         n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
         n2351, n2352, n2353, n2356, n2357, n2358, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2530, n2532, n2533, n2534, n2535, n2536,
         n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
         n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
         n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2703, n2705, n2707, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2777,
         n2778, n2779, n2780, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3,
         SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5,
         SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7,
         SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9,
         SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11,
         SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13,
         SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15,
         SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17,
         SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19,
         SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21,
         SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23,
         SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25,
         SYNOPSYS_UNCONNECTED_26, SYNOPSYS_UNCONNECTED_27, \shifter_0/n33 ,
         \shifter_0/n32 , \shifter_0/n31 , \shifter_0/n30 ,
         \shifter_0/o_shifted[4] , \shifter_0/n20 , \shifter_0/n19 ,
         \shifter_0/n18 , \shifter_0/n17 , \shifter_0/n16 , \shifter_0/n14 ,
         \shifter_0/n13 , \shifter_0/n12 , \shifter_0/n11 , \shifter_0/n10 ,
         \shifter_0/n9 , \shifter_0/n8 , \shifter_0/n7 , \shifter_0/n6 ,
         \shifter_0/n4 , \shifter_0/n1 , \shifter_0/n25 , \shifter_0/n24 ,
         \shifter_0/n21 , \shifter_0/shift_1b_0/n69 ,
         \shifter_0/shift_1b_0/n68 , \shifter_0/shift_1b_0/n67 ,
         \shifter_0/shift_1b_0/n66 , \shifter_0/shift_1b_0/n65 ,
         \shifter_0/shift_1b_0/n64 , \shifter_0/shift_1b_0/n63 ,
         \shifter_0/shift_1b_0/n62 , \shifter_0/shift_1b_0/n61 ,
         \shifter_0/shift_1b_0/n60 , \shifter_0/shift_1b_0/n59 ,
         \shifter_0/shift_1b_0/n58 , \shifter_0/shift_1b_0/n57 ,
         \shifter_0/shift_1b_0/n56 , \shifter_0/shift_1b_0/n55 ,
         \shifter_0/shift_1b_0/n54 , \shifter_0/shift_1b_0/n53 ,
         \shifter_0/shift_1b_0/n52 , \shifter_0/shift_1b_0/n51 ,
         \shifter_0/shift_1b_0/n50 , \shifter_0/shift_1b_0/n49 ,
         \shifter_0/shift_1b_0/n48 , \shifter_0/shift_1b_0/n47 ,
         \shifter_0/shift_1b_0/n46 , \shifter_0/shift_1b_0/n45 ,
         \shifter_0/shift_1b_0/n44 , \shifter_0/shift_1b_0/n43 ,
         \shifter_0/shift_1b_0/n42 , \shifter_0/shift_1b_0/n41 ,
         \shifter_0/shift_1b_0/n40 , \shifter_0/shift_1b_0/n39 ,
         \shifter_0/shift_1b_0/n38 , \shifter_0/shift_1b_0/n37 ,
         \shifter_0/shift_1b_0/n36 , \shifter_0/shift_1b_0/n35 ,
         \shifter_0/shift_1b_0/n34 , \shifter_0/shift_1b_0/n33 ,
         \shifter_0/shift_3b_0/n72 , \shifter_0/shift_3b_0/n71 ,
         \shifter_0/shift_3b_0/n70 , \shifter_0/shift_3b_0/n69 ,
         \shifter_0/shift_3b_0/n68 , \shifter_0/shift_3b_0/n67 ,
         \shifter_0/shift_3b_0/n66 , \shifter_0/shift_3b_0/n59 ,
         \shifter_0/shift_3b_0/n58 , \shifter_0/shift_3b_0/n57 ,
         \shifter_0/shift_3b_0/n56 , \shifter_0/shift_3b_0/n55 ,
         \shifter_0/shift_3b_0/n54 , \shifter_0/shift_3b_0/n53 ,
         \shifter_0/shift_3b_0/n52 , \shifter_0/shift_3b_0/n51 ,
         \shifter_0/shift_3b_0/n50 , \shifter_0/shift_3b_0/n49 ,
         \shifter_0/shift_3b_0/n48 , \shifter_0/shift_3b_0/n47 ,
         \shifter_0/shift_3b_0/n46 , \shifter_0/shift_3b_0/n45 ,
         \shifter_0/shift_3b_0/n44 , \shifter_0/shift_3b_0/n43 ,
         \shifter_0/shift_3b_0/n42 , \shifter_0/shift_3b_0/n41 ,
         \shifter_0/shift_3b_0/n40 , \shifter_0/shift_3b_0/n39 ,
         \shifter_0/shift_3b_0/n38 , \shifter_0/shift_3b_0/n37 ,
         \shifter_0/shift_3b_0/n36 , \shifter_0/shift_3b_0/n35 ,
         \shifter_0/shift_3b_0/n65 , \shifter_0/shift_3b_0/n64 ,
         \shifter_0/shift_3b_0/n63 , \shifter_0/shift_3b_0/n62 ,
         \shifter_0/shift_3b_0/n61 , \shifter_0/shift_3b_0/n60 ,
         \shifter_0/shift_3b_0/n13 , \shifter_0/shift_3b_0/n5 ,
         \shifter_0/shift_3b_0/n4 , \shifter_0/shift_3b_0/n3 ,
         \shifter_0/shift_3b_0/n2 , \shifter_0/shift_3b_0/n34 ,
         \shifter_0/shift_3b_0/n33 , \shifter_0/shift_3b_0/n32 ,
         \shifter_0/shift_3b_0/n31 , \shifter_0/shift_3b_0/n30 ,
         \shifter_0/shift_3b_0/n29 , \shifter_0/shift_3b_0/n28 ,
         \shifter_0/shift_3b_0/n27 , \shifter_0/shift_3b_0/n26 ,
         \shifter_0/shift_3b_0/n25 , \shifter_0/shift_3b_0/n24 ,
         \shifter_0/shift_3b_0/n23 , \shifter_0/shift_3b_0/n22 ,
         \shifter_0/shift_3b_0/n21 , \shifter_0/shift_3b_0/n20 ,
         \shifter_0/shift_3b_0/n19 , \shifter_0/shift_3b_0/n18 ,
         \shifter_0/shift_3b_0/n14 , \shifter_0/shift_3b_0/n12 ,
         \shifter_0/shift_3b_0/n11 , \shifter_0/shift_3b_0/n10 ,
         \shifter_0/shift_3b_0/n9 , \shifter_0/shift_3b_0/n8 ,
         \shifter_0/shift_3b_0/n7 , \shifter_0/shift_3b_0/n6 ,
         \shifter_0/shift_3b_0/shift1 , \shifter_0/shift_3b_0/shift_1b_0/n67 ,
         \shifter_0/shift_3b_0/shift_1b_0/n66 ,
         \shifter_0/shift_3b_0/shift_1b_0/n65 ,
         \shifter_0/shift_3b_0/shift_1b_0/n64 ,
         \shifter_0/shift_3b_0/shift_1b_0/n63 ,
         \shifter_0/shift_3b_0/shift_1b_0/n62 ,
         \shifter_0/shift_3b_0/shift_1b_0/n61 ,
         \shifter_0/shift_3b_0/shift_1b_0/n60 ,
         \shifter_0/shift_3b_0/shift_1b_0/n59 ,
         \shifter_0/shift_3b_0/shift_1b_0/n58 ,
         \shifter_0/shift_3b_0/shift_1b_0/n57 ,
         \shifter_0/shift_3b_0/shift_1b_0/n56 ,
         \shifter_0/shift_3b_0/shift_1b_0/n55 ,
         \shifter_0/shift_3b_0/shift_1b_0/n54 ,
         \shifter_0/shift_3b_0/shift_1b_0/n53 ,
         \shifter_0/shift_3b_0/shift_1b_0/n52 ,
         \shifter_0/shift_3b_0/shift_1b_0/n51 ,
         \shifter_0/shift_3b_0/shift_1b_0/n50 ,
         \shifter_0/shift_3b_0/shift_1b_0/n49 ,
         \shifter_0/shift_3b_0/shift_1b_0/n48 ,
         \shifter_0/shift_3b_0/shift_1b_0/n47 ,
         \shifter_0/shift_3b_0/shift_1b_0/n46 ,
         \shifter_0/shift_3b_0/shift_1b_0/n45 ,
         \shifter_0/shift_3b_0/shift_1b_0/n44 ,
         \shifter_0/shift_3b_0/shift_1b_0/n43 ,
         \shifter_0/shift_3b_0/shift_1b_0/n42 ,
         \shifter_0/shift_3b_0/shift_1b_0/n41 ,
         \shifter_0/shift_3b_0/shift_1b_0/n40 ,
         \shifter_0/shift_3b_0/shift_1b_0/n39 ,
         \shifter_0/shift_3b_0/shift_1b_0/n38 ,
         \shifter_0/shift_3b_0/shift_1b_0/n37 ,
         \shifter_0/shift_3b_0/shift_1b_0/n36 ,
         \shifter_0/shift_3b_0/shift_1b_0/n35 ,
         \shifter_0/shift_3b_0/shift_1b_0/n34 ,
         \shifter_0/shift_3b_0/shift_1b_0/n33 , \shifter_0/shift_3b_1/n72 ,
         \shifter_0/shift_3b_1/n71 , \shifter_0/shift_3b_1/n70 ,
         \shifter_0/shift_3b_1/n69 , \shifter_0/shift_3b_1/n68 ,
         \shifter_0/shift_3b_1/n67 , \shifter_0/shift_3b_1/n66 ,
         \shifter_0/shift_3b_1/n60 , \shifter_0/shift_3b_1/n59 ,
         \shifter_0/shift_3b_1/n58 , \shifter_0/shift_3b_1/n57 ,
         \shifter_0/shift_3b_1/n56 , \shifter_0/shift_3b_1/n55 ,
         \shifter_0/shift_3b_1/n54 , \shifter_0/shift_3b_1/n53 ,
         \shifter_0/shift_3b_1/n52 , \shifter_0/shift_3b_1/n51 ,
         \shifter_0/shift_3b_1/n50 , \shifter_0/shift_3b_1/n49 ,
         \shifter_0/shift_3b_1/n48 , \shifter_0/shift_3b_1/n47 ,
         \shifter_0/shift_3b_1/n46 , \shifter_0/shift_3b_1/n45 ,
         \shifter_0/shift_3b_1/n44 , \shifter_0/shift_3b_1/n43 ,
         \shifter_0/shift_3b_1/n42 , \shifter_0/shift_3b_1/n41 ,
         \shifter_0/shift_3b_1/n40 , \shifter_0/shift_3b_1/n39 ,
         \shifter_0/shift_3b_1/n38 , \shifter_0/shift_3b_1/n37 ,
         \shifter_0/shift_3b_1/n36 , \shifter_0/shift_3b_1/n35 ,
         \shifter_0/shift_3b_1/n65 , \shifter_0/shift_3b_1/n64 ,
         \shifter_0/shift_3b_1/n63 , \shifter_0/shift_3b_1/n62 ,
         \shifter_0/shift_3b_1/n61 , \shifter_0/shift_3b_1/n14 ,
         \shifter_0/shift_3b_1/n4 , \shifter_0/shift_3b_1/n3 ,
         \shifter_0/shift_3b_1/n2 , \shifter_0/shift_3b_1/n34 ,
         \shifter_0/shift_3b_1/n33 , \shifter_0/shift_3b_1/n32 ,
         \shifter_0/shift_3b_1/n31 , \shifter_0/shift_3b_1/n30 ,
         \shifter_0/shift_3b_1/n29 , \shifter_0/shift_3b_1/n28 ,
         \shifter_0/shift_3b_1/n27 , \shifter_0/shift_3b_1/n26 ,
         \shifter_0/shift_3b_1/n25 , \shifter_0/shift_3b_1/n24 ,
         \shifter_0/shift_3b_1/n23 , \shifter_0/shift_3b_1/n22 ,
         \shifter_0/shift_3b_1/n21 , \shifter_0/shift_3b_1/n20 ,
         \shifter_0/shift_3b_1/n19 , \shifter_0/shift_3b_1/n16 ,
         \shifter_0/shift_3b_1/n13 , \shifter_0/shift_3b_1/n12 ,
         \shifter_0/shift_3b_1/n11 , \shifter_0/shift_3b_1/n10 ,
         \shifter_0/shift_3b_1/n9 , \shifter_0/shift_3b_1/n8 ,
         \shifter_0/shift_3b_1/n7 , \shifter_0/shift_3b_1/n6 ,
         \shifter_0/shift_3b_1/n5 , \shifter_0/shift_3b_1/shift1 ,
         \shifter_0/shift_3b_1/shift_1b_0/n99 ,
         \shifter_0/shift_3b_1/shift_1b_0/n98 ,
         \shifter_0/shift_3b_1/shift_1b_0/n97 ,
         \shifter_0/shift_3b_1/shift_1b_0/n96 ,
         \shifter_0/shift_3b_1/shift_1b_0/n95 ,
         \shifter_0/shift_3b_1/shift_1b_0/n94 ,
         \shifter_0/shift_3b_1/shift_1b_0/n93 ,
         \shifter_0/shift_3b_1/shift_1b_0/n92 ,
         \shifter_0/shift_3b_1/shift_1b_0/n91 ,
         \shifter_0/shift_3b_1/shift_1b_0/n90 ,
         \shifter_0/shift_3b_1/shift_1b_0/n89 ,
         \shifter_0/shift_3b_1/shift_1b_0/n88 ,
         \shifter_0/shift_3b_1/shift_1b_0/n87 ,
         \shifter_0/shift_3b_1/shift_1b_0/n86 ,
         \shifter_0/shift_3b_1/shift_1b_0/n85 ,
         \shifter_0/shift_3b_1/shift_1b_0/n84 ,
         \shifter_0/shift_3b_1/shift_1b_0/n83 ,
         \shifter_0/shift_3b_1/shift_1b_0/n82 ,
         \shifter_0/shift_3b_1/shift_1b_0/n81 ,
         \shifter_0/shift_3b_1/shift_1b_0/n80 ,
         \shifter_0/shift_3b_1/shift_1b_0/n79 ,
         \shifter_0/shift_3b_1/shift_1b_0/n78 ,
         \shifter_0/shift_3b_1/shift_1b_0/n77 ,
         \shifter_0/shift_3b_1/shift_1b_0/n76 ,
         \shifter_0/shift_3b_1/shift_1b_0/n75 ,
         \shifter_0/shift_3b_1/shift_1b_0/n74 ,
         \shifter_0/shift_3b_1/shift_1b_0/n73 ,
         \shifter_0/shift_3b_1/shift_1b_0/n72 ,
         \shifter_0/shift_3b_1/shift_1b_0/n71 ,
         \shifter_0/shift_3b_1/shift_1b_0/n70 ,
         \shifter_0/shift_3b_1/shift_1b_0/n69 ,
         \shifter_0/shift_3b_1/shift_1b_0/n68 ,
         \shifter_0/shift_3b_1/shift_1b_0/n67 ,
         \shifter_0/shift_3b_1/shift_1b_0/n66 ,
         \shifter_0/shift_3b_1/shift_1b_0/n65 ,
         \shifter_0/shift_3b_1/shift_1b_0/n64 , \shifter_0/shift_7b_0/n80 ,
         \shifter_0/shift_7b_0/n79 , \shifter_0/shift_7b_0/n78 ,
         \shifter_0/shift_7b_0/n77 , \shifter_0/shift_7b_0/n76 ,
         \shifter_0/shift_7b_0/n75 , \shifter_0/shift_7b_0/n74 ,
         \shifter_0/shift_7b_0/n73 , \shifter_0/shift_7b_0/n72 ,
         \shifter_0/shift_7b_0/n71 , \shifter_0/shift_7b_0/n70 ,
         \shifter_0/shift_7b_0/n69 , \shifter_0/shift_7b_0/n68 ,
         \shifter_0/shift_7b_0/n56 , \shifter_0/shift_7b_0/n55 ,
         \shifter_0/shift_7b_0/n54 , \shifter_0/shift_7b_0/n53 ,
         \shifter_0/shift_7b_0/n52 , \shifter_0/shift_7b_0/n51 ,
         \shifter_0/shift_7b_0/n50 , \shifter_0/shift_7b_0/n49 ,
         \shifter_0/shift_7b_0/n48 , \shifter_0/shift_7b_0/n47 ,
         \shifter_0/shift_7b_0/n46 , \shifter_0/shift_7b_0/n45 ,
         \shifter_0/shift_7b_0/n44 , \shifter_0/shift_7b_0/n43 ,
         \shifter_0/shift_7b_0/n42 , \shifter_0/shift_7b_0/n41 ,
         \shifter_0/shift_7b_0/n40 , \shifter_0/shift_7b_0/n39 ,
         \shifter_0/shift_7b_0/n67 , \shifter_0/shift_7b_0/n66 ,
         \shifter_0/shift_7b_0/n65 , \shifter_0/shift_7b_0/n64 ,
         \shifter_0/shift_7b_0/n63 , \shifter_0/shift_7b_0/n62 ,
         \shifter_0/shift_7b_0/n61 , \shifter_0/shift_7b_0/n60 ,
         \shifter_0/shift_7b_0/n59 , \shifter_0/shift_7b_0/n58 ,
         \shifter_0/shift_7b_0/n57 , \shifter_0/shift_7b_0/n21 ,
         \shifter_0/shift_7b_0/n10 , \shifter_0/shift_7b_0/n9 ,
         \shifter_0/shift_7b_0/n8 , \shifter_0/shift_7b_0/n7 ,
         \shifter_0/shift_7b_0/n6 , \shifter_0/shift_7b_0/n5 ,
         \shifter_0/shift_7b_0/n4 , \shifter_0/shift_7b_0/n38 ,
         \shifter_0/shift_7b_0/n37 , \shifter_0/shift_7b_0/n36 ,
         \shifter_0/shift_7b_0/n35 , \shifter_0/shift_7b_0/n34 ,
         \shifter_0/shift_7b_0/n33 , \shifter_0/shift_7b_0/n32 ,
         \shifter_0/shift_7b_0/n31 , \shifter_0/shift_7b_0/n30 ,
         \shifter_0/shift_7b_0/n29 , \shifter_0/shift_7b_0/n20 ,
         \shifter_0/shift_7b_0/n19 , \shifter_0/shift_7b_0/n18 ,
         \shifter_0/shift_7b_0/n17 , \shifter_0/shift_7b_0/n16 ,
         \shifter_0/shift_7b_0/n15 , \shifter_0/shift_7b_0/n14 ,
         \shifter_0/shift_7b_0/n13 , \shifter_0/shift_7b_0/n12 ,
         \shifter_0/shift_7b_0/n11 , \shifter_0/shift_7b_0/shift_3b_0/n72 ,
         \shifter_0/shift_7b_0/shift_3b_0/n71 ,
         \shifter_0/shift_7b_0/shift_3b_0/n70 ,
         \shifter_0/shift_7b_0/shift_3b_0/n69 ,
         \shifter_0/shift_7b_0/shift_3b_0/n68 ,
         \shifter_0/shift_7b_0/shift_3b_0/n67 ,
         \shifter_0/shift_7b_0/shift_3b_0/n66 ,
         \shifter_0/shift_7b_0/shift_3b_0/n60 ,
         \shifter_0/shift_7b_0/shift_3b_0/n59 ,
         \shifter_0/shift_7b_0/shift_3b_0/n58 ,
         \shifter_0/shift_7b_0/shift_3b_0/n57 ,
         \shifter_0/shift_7b_0/shift_3b_0/n56 ,
         \shifter_0/shift_7b_0/shift_3b_0/n55 ,
         \shifter_0/shift_7b_0/shift_3b_0/n54 ,
         \shifter_0/shift_7b_0/shift_3b_0/n53 ,
         \shifter_0/shift_7b_0/shift_3b_0/n52 ,
         \shifter_0/shift_7b_0/shift_3b_0/n51 ,
         \shifter_0/shift_7b_0/shift_3b_0/n50 ,
         \shifter_0/shift_7b_0/shift_3b_0/n49 ,
         \shifter_0/shift_7b_0/shift_3b_0/n48 ,
         \shifter_0/shift_7b_0/shift_3b_0/n47 ,
         \shifter_0/shift_7b_0/shift_3b_0/n46 ,
         \shifter_0/shift_7b_0/shift_3b_0/n45 ,
         \shifter_0/shift_7b_0/shift_3b_0/n44 ,
         \shifter_0/shift_7b_0/shift_3b_0/n43 ,
         \shifter_0/shift_7b_0/shift_3b_0/n42 ,
         \shifter_0/shift_7b_0/shift_3b_0/n41 ,
         \shifter_0/shift_7b_0/shift_3b_0/n40 ,
         \shifter_0/shift_7b_0/shift_3b_0/n39 ,
         \shifter_0/shift_7b_0/shift_3b_0/n38 ,
         \shifter_0/shift_7b_0/shift_3b_0/n37 ,
         \shifter_0/shift_7b_0/shift_3b_0/n36 ,
         \shifter_0/shift_7b_0/shift_3b_0/n35 ,
         \shifter_0/shift_7b_0/shift_3b_0/n65 ,
         \shifter_0/shift_7b_0/shift_3b_0/n64 ,
         \shifter_0/shift_7b_0/shift_3b_0/n63 ,
         \shifter_0/shift_7b_0/shift_3b_0/n62 ,
         \shifter_0/shift_7b_0/shift_3b_0/n61 ,
         \shifter_0/shift_7b_0/shift_3b_0/n18 ,
         \shifter_0/shift_7b_0/shift_3b_0/n4 ,
         \shifter_0/shift_7b_0/shift_3b_0/n3 ,
         \shifter_0/shift_7b_0/shift_3b_0/n2 ,
         \shifter_0/shift_7b_0/shift_3b_0/n34 ,
         \shifter_0/shift_7b_0/shift_3b_0/n33 ,
         \shifter_0/shift_7b_0/shift_3b_0/n32 ,
         \shifter_0/shift_7b_0/shift_3b_0/n31 ,
         \shifter_0/shift_7b_0/shift_3b_0/n30 ,
         \shifter_0/shift_7b_0/shift_3b_0/n29 ,
         \shifter_0/shift_7b_0/shift_3b_0/n28 ,
         \shifter_0/shift_7b_0/shift_3b_0/n27 ,
         \shifter_0/shift_7b_0/shift_3b_0/n26 ,
         \shifter_0/shift_7b_0/shift_3b_0/n25 ,
         \shifter_0/shift_7b_0/shift_3b_0/n24 ,
         \shifter_0/shift_7b_0/shift_3b_0/n23 ,
         \shifter_0/shift_7b_0/shift_3b_0/n20 ,
         \shifter_0/shift_7b_0/shift_3b_0/n17 ,
         \shifter_0/shift_7b_0/shift_3b_0/n16 ,
         \shifter_0/shift_7b_0/shift_3b_0/n15 ,
         \shifter_0/shift_7b_0/shift_3b_0/n14 ,
         \shifter_0/shift_7b_0/shift_3b_0/n13 ,
         \shifter_0/shift_7b_0/shift_3b_0/n12 ,
         \shifter_0/shift_7b_0/shift_3b_0/n11 ,
         \shifter_0/shift_7b_0/shift_3b_0/n10 ,
         \shifter_0/shift_7b_0/shift_3b_0/n9 ,
         \shifter_0/shift_7b_0/shift_3b_0/n8 ,
         \shifter_0/shift_7b_0/shift_3b_0/n7 ,
         \shifter_0/shift_7b_0/shift_3b_0/n6 ,
         \shifter_0/shift_7b_0/shift_3b_0/n5 ,
         \shifter_0/shift_7b_0/shift_3b_0/shift1 ,
         \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n67 ,
         \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n66 ,
         \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n65 ,
         \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n64 ,
         \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n63 ,
         \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n62 ,
         \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n61 ,
         \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n60 ,
         \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n59 ,
         \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n58 ,
         \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n57 ,
         \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n56 ,
         \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n55 ,
         \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n54 ,
         \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n53 ,
         \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n52 ,
         \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n51 ,
         \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n50 ,
         \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n49 ,
         \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n48 ,
         \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n47 ,
         \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n46 ,
         \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n45 ,
         \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n44 ,
         \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n43 ,
         \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n42 ,
         \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n41 ,
         \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n40 ,
         \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n39 ,
         \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n38 ,
         \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n37 ,
         \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n36 ,
         \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n35 ,
         \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n34 ,
         \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n33 , \adder_0/G6_1 ,
         \adder_0/G6_3 , \adder_0/G6_5 , \adder_0/G6_7 , \adder_0/G6_9 ,
         \adder_0/G6_11 , \adder_0/G6_13 , \adder_0/G6_15 , \adder_0/G6_17 ,
         \adder_0/G6_19 , \adder_0/G6_21 , \adder_0/G6_23 , \adder_0/G6_25 ,
         \adder_0/G6_27 , \adder_0/G6_29_ , \adder_0/G5[8] , \adder_0/G5[9] ,
         \adder_0/G5[10] , \adder_0/G5[11] , \adder_0/G5[12] ,
         \adder_0/G5[13] , \adder_0/G5[14] , \adder_0/G5[15] , \adder_0/G4[4] ,
         \adder_0/G4[5] , \adder_0/G4[6] , \adder_0/G4[7] , \adder_0/G4[8] ,
         \adder_0/G4[9] , \adder_0/G4[10] , \adder_0/G4[11] , \adder_0/G4[12] ,
         \adder_0/G4[13] , \adder_0/G4[14] , \adder_0/G4[15] , \adder_0/P3[4] ,
         \adder_0/P3[5] , \adder_0/P3[6] , \adder_0/P3[7] , \adder_0/P3[8] ,
         \adder_0/P3[9] , \adder_0/P3[10] , \adder_0/P3[11] , \adder_0/P3[12] ,
         \adder_0/P3[13] , \adder_0/P3[14] , \adder_0/P3[15] , \adder_0/G3[2] ,
         \adder_0/G3[3] , \adder_0/G3[4] , \adder_0/G3[5] , \adder_0/G3[6] ,
         \adder_0/G3[7] , \adder_0/G3[8] , \adder_0/G3[9] , \adder_0/G3[10] ,
         \adder_0/G3[11] , \adder_0/G3[12] , \adder_0/G3[13] ,
         \adder_0/G3[14] , \adder_0/G3[15] , \adder_0/P2[2] , \adder_0/P2[3] ,
         \adder_0/P2[4] , \adder_0/P2[5] , \adder_0/P2[6] , \adder_0/P2[7] ,
         \adder_0/P2[8] , \adder_0/P2[9] , \adder_0/P2[10] , \adder_0/P2[11] ,
         \adder_0/P2[12] , \adder_0/P2[13] , \adder_0/P2[14] ,
         \adder_0/P2[15] , \adder_0/G2[1] , \adder_0/G2[2] , \adder_0/G2[3] ,
         \adder_0/G2[4] , \adder_0/G2[5] , \adder_0/G2[6] , \adder_0/G2[7] ,
         \adder_0/G2[8] , \adder_0/G2[9] , \adder_0/G2[10] , \adder_0/G2[11] ,
         \adder_0/G2[12] , \adder_0/G2[13] , \adder_0/G2[14] ,
         \adder_0/G2[15] , \adder_0/P1[1] , \adder_0/P1[2] , \adder_0/P1[3] ,
         \adder_0/P1[4] , \adder_0/P1[5] , \adder_0/P1[6] , \adder_0/P1[7] ,
         \adder_0/P1[8] , \adder_0/P1[9] , \adder_0/P1[10] , \adder_0/P1[11] ,
         \adder_0/P1[12] , \adder_0/P1[13] , \adder_0/P1[14] ,
         \adder_0/P1[15] , \adder_0/G1[0] , \adder_0/G1[1] , \adder_0/G1[2] ,
         \adder_0/G1[3] , \adder_0/G1[4] , \adder_0/G1[5] , \adder_0/G1[6] ,
         \adder_0/G1[7] , \adder_0/G1[8] , \adder_0/G1[9] , \adder_0/G1[10] ,
         \adder_0/G1[11] , \adder_0/G1[12] , \adder_0/G1[13] ,
         \adder_0/G1[14] , \adder_0/G1[15] , \adder_0/G0[0] , \adder_0/G0[1] ,
         \adder_0/G0[2] , \adder_0/G0[3] , \adder_0/G0[4] , \adder_0/G0[5] ,
         \adder_0/G0[6] , \adder_0/G0[7] , \adder_0/G0[8] , \adder_0/G0[9] ,
         \adder_0/G0[10] , \adder_0/G0[11] , \adder_0/G0[12] ,
         \adder_0/G0[13] , \adder_0/G0[14] , \adder_0/G0[15] ,
         \adder_0/G0[16] , \adder_0/G0[17] , \adder_0/G0[18] ,
         \adder_0/G0[19] , \adder_0/G0[20] , \adder_0/G0[21] ,
         \adder_0/G0[22] , \adder_0/G0[23] , \adder_0/G0[24] ,
         \adder_0/G0[25] , \adder_0/G0[26] , \adder_0/G0[27] ,
         \adder_0/G0[28] , \adder_0/G0[29] , \adder_0/G0[30] ,
         \adder_0/G0[31] , \adder_0/P0[0] , \adder_0/P0[1] , \adder_0/P0[2] ,
         \adder_0/P0[3] , \adder_0/P0[4] , \adder_0/P0[5] , \adder_0/P0[6] ,
         \adder_0/P0[7] , \adder_0/P0[8] , \adder_0/P0[9] , \adder_0/P0[10] ,
         \adder_0/P0[11] , \adder_0/P0[12] , \adder_0/P0[13] ,
         \adder_0/P0[14] , \adder_0/P0[15] , \adder_0/P0[16] ,
         \adder_0/P0[17] , \adder_0/P0[18] , \adder_0/P0[19] ,
         \adder_0/P0[20] , \adder_0/P0[21] , \adder_0/P0[22] ,
         \adder_0/P0[23] , \adder_0/P0[24] , \adder_0/P0[25] ,
         \adder_0/P0[26] , \adder_0/P0[27] , \adder_0/P0[28] ,
         \adder_0/P0[29] , \adder_0/P0[30] , \adder_0/P0[31] , \adder_0/o_c ,
         \adder_0/operator_C_stage_1_0/n2 , \adder_0/operator_B_stage_1_1/n2 ,
         \adder_0/operator_B_stage_1_2/n3 , \adder_0/operator_B_stage_1_3/n3 ,
         \adder_0/operator_B_stage_1_4/n3 , \adder_0/operator_B_stage_1_5/n3 ,
         \adder_0/operator_B_stage_1_6/n3 , \adder_0/operator_B_stage_1_7/n3 ,
         \adder_0/operator_B_stage_1_8/n3 , \adder_0/operator_B_stage_1_9/n3 ,
         \adder_0/operator_B_stage_1_10/n3 ,
         \adder_0/operator_B_stage_1_11/n3 ,
         \adder_0/operator_B_stage_1_12/n3 ,
         \adder_0/operator_B_stage_1_13/n3 ,
         \adder_0/operator_B_stage_1_14/n3 ,
         \adder_0/operator_B_stage_1_15/n3 , \adder_0/operator_C_stage_2_1/n3 ,
         \adder_0/operator_B_stage_2_2/n3 , \adder_0/operator_B_stage_2_3/n3 ,
         \adder_0/operator_B_stage_2_4/n3 , \adder_0/operator_B_stage_2_5/n3 ,
         \adder_0/operator_B_stage_2_6/n3 , \adder_0/operator_B_stage_2_7/n3 ,
         \adder_0/operator_B_stage_2_8/n3 , \adder_0/operator_B_stage_2_9/n3 ,
         \adder_0/operator_B_stage_2_10/n3 ,
         \adder_0/operator_B_stage_2_11/n3 ,
         \adder_0/operator_B_stage_2_12/n3 ,
         \adder_0/operator_B_stage_2_13/n3 ,
         \adder_0/operator_B_stage_2_14/n3 ,
         \adder_0/operator_B_stage_2_15/n3 , \adder_0/operator_C_stage_3_2/n3 ,
         \adder_0/operator_C_stage_3_3/n3 , \adder_0/operator_B_stage_3_4/n3 ,
         \adder_0/operator_B_stage_3_5/n3 , \adder_0/operator_B_stage_3_6/n3 ,
         \adder_0/operator_B_stage_3_7/n3 , \adder_0/operator_B_stage_3_8/n3 ,
         \adder_0/operator_B_stage_3_9/n3 , \adder_0/operator_B_stage_3_10/n3 ,
         \adder_0/operator_B_stage_3_11/n3 ,
         \adder_0/operator_B_stage_3_12/n3 ,
         \adder_0/operator_B_stage_3_13/n3 ,
         \adder_0/operator_B_stage_3_14/n3 ,
         \adder_0/operator_B_stage_3_15/n3 , \adder_0/operator_C_stage_4_4/n3 ,
         \adder_0/operator_C_stage_4_5/n3 , \adder_0/operator_C_stage_4_6/n3 ,
         \adder_0/operator_C_stage_4_7/n3 , \adder_0/operator_B_stage_4_8/n3 ,
         \adder_0/operator_B_stage_4_9/n3 , \adder_0/operator_B_stage_4_10/n3 ,
         \adder_0/operator_B_stage_4_11/n3 ,
         \adder_0/operator_B_stage_4_12/n3 ,
         \adder_0/operator_B_stage_4_13/n3 ,
         \adder_0/operator_B_stage_4_14/n3 ,
         \adder_0/operator_B_stage_4_15/n3 , \adder_0/operator_C_stage_5_8/n3 ,
         \adder_0/operator_C_stage_5_9/n3 , \adder_0/operator_C_stage_5_10/n3 ,
         \adder_0/operator_C_stage_5_11/n3 ,
         \adder_0/operator_C_stage_5_12/n3 ,
         \adder_0/operator_C_stage_5_13/n3 ,
         \adder_0/operator_C_stage_5_14/n3 ,
         \adder_0/operator_C_stage_5_15/n3 , \adder_0/operator_C_stage_6_0/n3 ,
         \adder_0/operator_C_stage_6_1/n3 , \adder_0/operator_C_stage_6_2/n3 ,
         \adder_0/operator_C_stage_6_3/n3 , \adder_0/operator_C_stage_6_4/n3 ,
         \adder_0/operator_C_stage_6_5/n3 , \adder_0/operator_C_stage_6_6/n3 ,
         \adder_0/operator_C_stage_6_7/n3 , \adder_0/operator_C_stage_6_8/n3 ,
         \adder_0/operator_C_stage_6_9/n3 , \adder_0/operator_C_stage_6_10/n3 ,
         \adder_0/operator_C_stage_6_11/n3 ,
         \adder_0/operator_C_stage_6_12/n3 ,
         \adder_0/operator_C_stage_6_13/n3 ,
         \adder_0/operator_C_stage_6_14/n3 ,
         \adder_0/operator_C_stage_6_15/n3 , \adder_1/G6_1 , \adder_1/G6_3 ,
         \adder_1/G6_5 , \adder_1/G6_7 , \adder_1/G6_9 , \adder_1/G6_11 ,
         \adder_1/G6_13 , \adder_1/G6_15 , \adder_1/G6_17 , \adder_1/G6_19 ,
         \adder_1/G6_21 , \adder_1/G6_23 , \adder_1/G6_25 , \adder_1/G6_27 ,
         \adder_1/G6_29_ , \adder_1/G5[8] , \adder_1/G5[9] , \adder_1/G5[10] ,
         \adder_1/G5[11] , \adder_1/G5[12] , \adder_1/G5[13] ,
         \adder_1/G5[14] , \adder_1/G5[15] , \adder_1/G4[4] , \adder_1/G4[5] ,
         \adder_1/G4[6] , \adder_1/G4[7] , \adder_1/G4[8] , \adder_1/G4[9] ,
         \adder_1/G4[10] , \adder_1/G4[11] , \adder_1/G4[12] ,
         \adder_1/G4[13] , \adder_1/G4[14] , \adder_1/G4[15] , \adder_1/P3[4] ,
         \adder_1/P3[5] , \adder_1/P3[6] , \adder_1/P3[7] , \adder_1/P3[8] ,
         \adder_1/P3[9] , \adder_1/P3[10] , \adder_1/P3[11] , \adder_1/P3[12] ,
         \adder_1/P3[13] , \adder_1/P3[14] , \adder_1/P3[15] , \adder_1/G3[2] ,
         \adder_1/G3[3] , \adder_1/G3[4] , \adder_1/G3[5] , \adder_1/G3[6] ,
         \adder_1/G3[7] , \adder_1/G3[8] , \adder_1/G3[9] , \adder_1/G3[10] ,
         \adder_1/G3[11] , \adder_1/G3[12] , \adder_1/G3[13] ,
         \adder_1/G3[14] , \adder_1/G3[15] , \adder_1/P2[2] , \adder_1/P2[3] ,
         \adder_1/P2[4] , \adder_1/P2[5] , \adder_1/P2[6] , \adder_1/P2[7] ,
         \adder_1/P2[8] , \adder_1/P2[9] , \adder_1/P2[10] , \adder_1/P2[11] ,
         \adder_1/P2[12] , \adder_1/P2[13] , \adder_1/P2[14] ,
         \adder_1/P2[15] , \adder_1/G2[1] , \adder_1/G2[2] , \adder_1/G2[3] ,
         \adder_1/G2[4] , \adder_1/G2[5] , \adder_1/G2[6] , \adder_1/G2[7] ,
         \adder_1/G2[8] , \adder_1/G2[9] , \adder_1/G2[10] , \adder_1/G2[11] ,
         \adder_1/G2[12] , \adder_1/G2[13] , \adder_1/G2[14] ,
         \adder_1/G2[15] , \adder_1/P1[1] , \adder_1/P1[2] , \adder_1/P1[3] ,
         \adder_1/P1[4] , \adder_1/P1[5] , \adder_1/P1[6] , \adder_1/P1[7] ,
         \adder_1/P1[8] , \adder_1/P1[9] , \adder_1/P1[10] , \adder_1/P1[11] ,
         \adder_1/P1[12] , \adder_1/P1[13] , \adder_1/P1[14] ,
         \adder_1/P1[15] , \adder_1/G1[0] , \adder_1/G1[1] , \adder_1/G1[2] ,
         \adder_1/G1[3] , \adder_1/G1[4] , \adder_1/G1[5] , \adder_1/G1[6] ,
         \adder_1/G1[7] , \adder_1/G1[8] , \adder_1/G1[9] , \adder_1/G1[10] ,
         \adder_1/G1[11] , \adder_1/G1[12] , \adder_1/G1[13] ,
         \adder_1/G1[14] , \adder_1/G1[15] , \adder_1/G0[0] , \adder_1/G0[1] ,
         \adder_1/G0[2] , \adder_1/G0[3] , \adder_1/G0[4] , \adder_1/G0[5] ,
         \adder_1/G0[6] , \adder_1/G0[7] , \adder_1/G0[8] , \adder_1/G0[9] ,
         \adder_1/G0[10] , \adder_1/G0[11] , \adder_1/G0[12] ,
         \adder_1/G0[13] , \adder_1/G0[14] , \adder_1/G0[15] ,
         \adder_1/G0[16] , \adder_1/G0[17] , \adder_1/G0[18] ,
         \adder_1/G0[19] , \adder_1/G0[20] , \adder_1/G0[21] ,
         \adder_1/G0[22] , \adder_1/G0[23] , \adder_1/G0[24] ,
         \adder_1/G0[25] , \adder_1/G0[26] , \adder_1/G0[27] ,
         \adder_1/G0[28] , \adder_1/G0[29] , \adder_1/G0[30] ,
         \adder_1/G0[31] , \adder_1/P0[0] , \adder_1/P0[1] , \adder_1/P0[2] ,
         \adder_1/P0[3] , \adder_1/P0[4] , \adder_1/P0[5] , \adder_1/P0[6] ,
         \adder_1/P0[7] , \adder_1/P0[8] , \adder_1/P0[9] , \adder_1/P0[10] ,
         \adder_1/P0[11] , \adder_1/P0[12] , \adder_1/P0[13] ,
         \adder_1/P0[14] , \adder_1/P0[15] , \adder_1/P0[16] ,
         \adder_1/P0[17] , \adder_1/P0[18] , \adder_1/P0[19] ,
         \adder_1/P0[20] , \adder_1/P0[21] , \adder_1/P0[22] ,
         \adder_1/P0[23] , \adder_1/P0[24] , \adder_1/P0[25] ,
         \adder_1/P0[26] , \adder_1/P0[27] , \adder_1/P0[28] ,
         \adder_1/P0[29] , \adder_1/P0[30] , \adder_1/P0[31] , \adder_1/o_c ,
         \adder_1/operator_C_stage_1_0/n3 , \adder_1/operator_B_stage_1_1/n3 ,
         \adder_1/operator_B_stage_1_2/n3 , \adder_1/operator_B_stage_1_3/n3 ,
         \adder_1/operator_B_stage_1_4/n3 , \adder_1/operator_B_stage_1_5/n3 ,
         \adder_1/operator_B_stage_1_6/n3 , \adder_1/operator_B_stage_1_7/n3 ,
         \adder_1/operator_B_stage_1_8/n3 , \adder_1/operator_B_stage_1_9/n3 ,
         \adder_1/operator_B_stage_1_10/n3 ,
         \adder_1/operator_B_stage_1_11/n3 ,
         \adder_1/operator_B_stage_1_12/n3 ,
         \adder_1/operator_B_stage_1_13/n3 ,
         \adder_1/operator_B_stage_1_14/n3 ,
         \adder_1/operator_B_stage_1_15/n3 , \adder_1/operator_C_stage_2_1/n3 ,
         \adder_1/operator_B_stage_2_2/n3 , \adder_1/operator_B_stage_2_3/n3 ,
         \adder_1/operator_B_stage_2_4/n3 , \adder_1/operator_B_stage_2_5/n3 ,
         \adder_1/operator_B_stage_2_6/n3 , \adder_1/operator_B_stage_2_7/n3 ,
         \adder_1/operator_B_stage_2_8/n3 , \adder_1/operator_B_stage_2_9/n3 ,
         \adder_1/operator_B_stage_2_10/n3 ,
         \adder_1/operator_B_stage_2_11/n3 ,
         \adder_1/operator_B_stage_2_12/n3 ,
         \adder_1/operator_B_stage_2_13/n3 ,
         \adder_1/operator_B_stage_2_14/n3 ,
         \adder_1/operator_B_stage_2_15/n3 , \adder_1/operator_C_stage_3_2/n3 ,
         \adder_1/operator_C_stage_3_3/n3 , \adder_1/operator_B_stage_3_4/n3 ,
         \adder_1/operator_B_stage_3_5/n3 , \adder_1/operator_B_stage_3_6/n3 ,
         \adder_1/operator_B_stage_3_7/n3 , \adder_1/operator_B_stage_3_8/n3 ,
         \adder_1/operator_B_stage_3_9/n3 , \adder_1/operator_B_stage_3_10/n3 ,
         \adder_1/operator_B_stage_3_11/n3 ,
         \adder_1/operator_B_stage_3_12/n3 ,
         \adder_1/operator_B_stage_3_13/n3 ,
         \adder_1/operator_B_stage_3_14/n3 ,
         \adder_1/operator_B_stage_3_15/n3 , \adder_1/operator_C_stage_4_4/n3 ,
         \adder_1/operator_C_stage_4_5/n3 , \adder_1/operator_C_stage_4_6/n3 ,
         \adder_1/operator_C_stage_4_7/n3 , \adder_1/operator_B_stage_4_8/n3 ,
         \adder_1/operator_B_stage_4_9/n3 , \adder_1/operator_B_stage_4_10/n3 ,
         \adder_1/operator_B_stage_4_11/n3 ,
         \adder_1/operator_B_stage_4_12/n3 ,
         \adder_1/operator_B_stage_4_13/n3 ,
         \adder_1/operator_B_stage_4_14/n3 ,
         \adder_1/operator_B_stage_4_15/n3 , \adder_1/operator_C_stage_5_8/n3 ,
         \adder_1/operator_C_stage_5_9/n3 , \adder_1/operator_C_stage_5_10/n3 ,
         \adder_1/operator_C_stage_5_11/n3 ,
         \adder_1/operator_C_stage_5_12/n3 ,
         \adder_1/operator_C_stage_5_13/n3 ,
         \adder_1/operator_C_stage_5_14/n3 ,
         \adder_1/operator_C_stage_5_15/n3 , \adder_1/operator_C_stage_6_0/n3 ,
         \adder_1/operator_C_stage_6_1/n3 , \adder_1/operator_C_stage_6_2/n3 ,
         \adder_1/operator_C_stage_6_3/n3 , \adder_1/operator_C_stage_6_4/n3 ,
         \adder_1/operator_C_stage_6_5/n3 , \adder_1/operator_C_stage_6_6/n3 ,
         \adder_1/operator_C_stage_6_7/n3 , \adder_1/operator_C_stage_6_8/n3 ,
         \adder_1/operator_C_stage_6_9/n3 , \adder_1/operator_C_stage_6_10/n3 ,
         \adder_1/operator_C_stage_6_11/n3 ,
         \adder_1/operator_C_stage_6_12/n3 ,
         \adder_1/operator_C_stage_6_13/n3 ,
         \adder_1/operator_C_stage_6_14/n3 ,
         \adder_1/operator_C_stage_6_15/n3 , \sra_198/n289 , \sra_198/n288 ,
         \sra_198/n287 , \sra_198/n286 , \sra_198/n285 , \sra_198/n284 ,
         \sra_198/n283 , \sra_198/n282 , \sra_198/n281 , \sra_198/n280 ,
         \sra_198/n279 , \sra_198/n278 , \sra_198/n277 , \sra_198/n276 ,
         \sra_198/n275 , \sra_198/n274 , \sra_198/n273 , \sra_198/n272 ,
         \sra_198/n271 , \sra_198/n270 , \sra_198/n269 , \sra_198/n268 ,
         \sra_198/n267 , \sra_198/n266 , \sra_198/n265 , \sra_198/n264 ,
         \sra_198/n263 , \sra_198/n262 , \sra_198/n261 , \sra_198/n260 ,
         \sra_198/n259 , \sra_198/n258 , \sra_198/n257 , \sra_198/n256 ,
         \sra_198/n255 , \sra_198/n254 , \sra_198/n253 , \sra_198/n252 ,
         \sra_198/n251 , \sra_198/n250 , \sra_198/n249 , \sra_198/n248 ,
         \sra_198/n247 , \sra_198/n246 , \sra_198/n245 , \sra_198/n244 ,
         \sra_198/n243 , \sra_198/n242 , \sra_198/n241 , \sra_198/n240 ,
         \sra_198/n239 , \sra_198/n238 , \sra_198/n237 , \sra_198/n236 ,
         \sra_198/n235 , \sra_198/n234 , \sra_198/n233 , \sra_198/n232 ,
         \sra_198/n231 , \sra_198/n230 , \sra_198/n229 , \sra_198/n228 ,
         \sra_198/n227 , \sra_198/n226 , \sra_198/n225 , \sra_198/n224 ,
         \sra_198/n223 , \sra_198/n222 , \sra_198/n221 , \sra_198/n220 ,
         \sra_198/n219 , \sra_198/n218 , \sra_198/n217 , \sra_198/n216 ,
         \sra_198/n215 , \sra_198/n214 , \sra_198/n212 , \sra_198/n211 ,
         \sra_198/n210 , \sra_198/n209 , \sra_198/n208 , \sra_198/n207 ,
         \sra_198/n206 , \sra_198/n205 , \sra_198/n204 , \sra_198/n203 ,
         \sra_198/n202 , \sra_198/n201 , \sra_198/n200 , \sra_198/n199 ,
         \sra_198/n198 , \sra_198/n197 , \sra_198/n196 , \sra_198/n195 ,
         \sra_198/n194 , \sra_198/n193 , \sra_198/n192 , \sra_198/n191 ,
         \sra_198/n190 , \sra_198/n189 , \sra_198/n188 , \sra_198/n187 ,
         \sra_198/n186 , \sra_198/n185 , \sra_198/n184 , \sra_198/n183 ,
         \sra_198/n182 , \sra_198/n181 , \sra_198/n180 , \sra_198/n179 ,
         \sra_198/n178 , \sra_198/n177 , \sra_198/n176 , \sra_198/n175 ,
         \sra_198/n174 , \sra_198/n173 , \sra_198/n172 , \sra_198/n171 ,
         \sra_198/n170 , \sra_198/n169 , \sra_198/n168 , \sra_198/n167 ,
         \sra_198/n166 , \sra_198/n165 , \sra_198/n164 , \sra_198/n163 ,
         \sra_198/n162 , \sra_198/n161 , \sra_198/n160 , \sra_198/n159 ,
         \sra_198/n158 , \sra_198/n157 , \sra_198/n156 , \sra_198/n155 ,
         \sra_198/n154 , \sra_198/n153 , \sra_198/n152 , \sra_198/n151 ,
         \sra_198/n150 , \sra_198/n149 , \sra_198/n148 , \sra_198/n147 ,
         \sra_198/n146 , \sra_198/n145 , \sra_198/n144 , \sra_198/n143 ,
         \sra_198/n142 , \sra_198/n141 , \sra_198/n140 , \sra_198/n139 ,
         \sra_198/n138 , \sra_198/n137 , \sra_198/n136 , \sra_198/n135 ,
         \sra_198/n134 , \sra_198/n133 , \sra_198/n132 , \sra_198/n131 ,
         \sra_198/n130 , \sra_198/n129 , \sra_198/n128 , \sra_198/n127 ,
         \sra_198/n126 , \sra_198/n125 , \sra_198/n124 , \sra_198/n123 ,
         \sra_198/n122 , \sra_198/n121 , \sra_198/n120 , \sra_198/n119 ,
         \sra_198/n118 , \sra_198/n117 , \sra_198/n116 , \sra_198/n115 ,
         \sra_198/n114 , \sra_198/n113 , \sra_198/n112 , \sra_198/n111 ,
         \sra_198/n110 , \sra_198/n109 , \sra_198/n108 , \sra_198/n107 ,
         \sra_198/n106 , \sra_198/n105 , \sra_198/n104 , \sra_198/n103 ,
         \sra_198/n102 , \sra_198/n101 , \sra_198/n100 , \sra_198/n99 ,
         \sra_198/n98 , \sra_198/n97 , \sra_198/n96 , \sra_198/n95 ,
         \sra_198/n94 , \sra_198/n93 , \sra_198/n92 , \sra_198/n91 ,
         \sra_198/n90 , \sra_198/n89 , \sra_198/n88 , \sra_198/n87 ,
         \sra_198/n86 , \sra_198/n85 , \sra_198/n84 , \sra_198/n83 ,
         \sra_198/n82 , \sra_198/n81 , \sra_198/n80 , \sra_198/n79 ,
         \sra_198/n78 , \sra_198/n77 , \sra_198/n76 , \sra_198/n75 ,
         \sra_198/n74 , \add_35/n3 , \add_35/n2 , \add_35/carry[3] ,
         \add_35/carry[4] , \add_35/carry[5] , \add_35/carry[6] ,
         \add_35/carry[7] , \add_35/carry[8] , \add_35/carry[9] ,
         \add_35/carry[10] , \add_35/carry[11] , \add_35/carry[12] ,
         \add_35/carry[13] , \add_35/carry[14] , \add_35/carry[15] ,
         \add_35/carry[16] , \add_35/carry[17] , \add_35/carry[18] ,
         \add_35/carry[19] , \add_35/carry[20] , \add_35/carry[21] ,
         \add_35/carry[22] , \add_35/carry[23] , \add_35/carry[24] ,
         \add_35/carry[25] , \add_35/carry[26] , \add_35/carry[27] ,
         \add_35/carry[28] , \add_35/carry[29] , \add_35/carry[30] ,
         \add_34/n6 , \add_34/n5 , \add_34/n4 , \add_34/n3 , \add_34/n2 ,
         \add_34/carry[3] , \add_34/carry[4] , \add_34/carry[5] ,
         \add_34/carry[6] , \add_34/carry[7] , \add_34/carry[8] ,
         \add_34/carry[9] , \add_34/carry[10] , \add_34/carry[11] ,
         \add_34/carry[12] , \add_34/carry[13] , \add_34/carry[14] ,
         \add_34/carry[15] , \add_34/carry[16] , \add_34/carry[17] ,
         \add_34/carry[18] , \add_34/carry[19] , \add_34/carry[20] ,
         \add_34/carry[21] , \add_34/carry[22] , \add_34/carry[23] ,
         \add_34/carry[24] , \add_34/carry[25] , \add_34/carry[26] ,
         \add_34/carry[27] , \add_34/carry[28] , \add_34/carry[29] ,
         \add_34/carry[30] ;
  wire   [30:2] nq;
  wire   [30:0] nqp1;
  wire   [30:0] q;
  wire   [30:0] qp1;
  wire   [31:0] sdata;
  wire   [31:0] sdata_o;
  wire   [3:0] shifted_o;
  wire   [5:0] state;
  wire   [5:0] ct_1;
  wire   [31:0] PR_1;
  wire   [31:0] reg_a;
  wire   [31:0] reg_b;
  wire   [31:0] sum;
  wire   [5:0] sum_ct;
  wire   [5:0] ct;
  wire   [31:0] \shifter_0/data_3 ;
  wire   [31:0] \shifter_0/data_2 ;
  wire   [31:0] \shifter_0/data_1 ;
  wire   [1:0] \shifter_0/shift_3b_0/data1 ;
  wire   [1:0] \shifter_0/shift_3b_1/data1 ;
  wire   [2:0] \shifter_0/shift_7b_0/shift1 ;
  wire   [3:0] \shifter_0/shift_7b_0/data1 ;
  wire   [1:0] \shifter_0/shift_7b_0/shift_3b_0/data1 ;
  wire   [15:8] \adder_0/P4 ;
  wire   [15:8] \adder_1/P4 ;

  SDFFR_X1 state_reg_reg_1_ ( .D(1'b1), .SI(n977), .SE(n941), .CK(i_clk), .RN(
        n3013), .Q(state_reg_1_0), .QN(n2929) );
  NAND3_X1 U2099 ( .A1(n935), .A2(n2320), .A3(n936), .ZN(n2489) );
  NAND3_X1 U2100 ( .A1(n2320), .A2(ct[3]), .A3(n935), .ZN(n2498) );
  NAND3_X1 U2101 ( .A1(n2320), .A2(ct[4]), .A3(n936), .ZN(n2499) );
  NAND3_X1 U2102 ( .A1(ct[1]), .A2(ct[0]), .A3(ct[2]), .ZN(n2497) );
  NAND3_X1 U2103 ( .A1(n938), .A2(n937), .A3(n939), .ZN(n2490) );
  NAND3_X1 U2104 ( .A1(n937), .A2(ct[0]), .A3(n938), .ZN(n2491) );
  NAND3_X1 U2105 ( .A1(n937), .A2(ct[1]), .A3(n939), .ZN(n2492) );
  NAND3_X1 U2106 ( .A1(ct[1]), .A2(ct[0]), .A3(n937), .ZN(n2493) );
  NAND3_X1 U2107 ( .A1(n938), .A2(ct[2]), .A3(n939), .ZN(n2494) );
  NAND3_X1 U2108 ( .A1(ct[2]), .A2(ct[0]), .A3(n938), .ZN(n2495) );
  NAND3_X1 U2109 ( .A1(ct[4]), .A2(ct[3]), .A3(n2320), .ZN(n2500) );
  NAND3_X1 U2110 ( .A1(ct[2]), .A2(ct[1]), .A3(n939), .ZN(n2496) );
  NAND3_X1 U2111 ( .A1(n2614), .A2(n2615), .A3(n3186), .ZN(n2610) );
  NAND3_X1 U2112 ( .A1(n2501), .A2(n2615), .A3(n2614), .ZN(n2401) );
  NAND3_X1 U2113 ( .A1(n2410), .A2(n2409), .A3(n3111), .ZN(n2344) );
  DFFS_X1 state_reg_0_ ( .D(n1191), .CK(i_clk), .SN(i_rst), .Q(state[0]), .QN(
        n3106) );
  DFFR_X1 DD_sign_reg ( .D(n1227), .CK(i_clk), .RN(n3000), .Q(), .QN(n2768) );
  DFFR_X1 ct_1_en_reg ( .D(n1113), .CK(i_clk), .RN(n3001), .Q(), .QN(n2769) );
  DFFR_X1 state_reg_reg_0_ ( .D(n1293), .CK(i_clk), .RN(n3000), .Q(), .QN(n941) );
  DFFR_X1 DR_reg_7_ ( .D(n1148), .CK(i_clk), .RN(n2995), .Q(n3138), .QN(n2713)
         );
  DFFR_X1 DR_reg_6_ ( .D(n1149), .CK(i_clk), .RN(n2994), .Q(n3136), .QN(n2712)
         );
  DFFR_X1 DR_reg_5_ ( .D(n1150), .CK(i_clk), .RN(n2992), .Q(n3134), .QN(n2711)
         );
  DFFR_X1 DR_reg_4_ ( .D(n1151), .CK(i_clk), .RN(n2986), .Q(n3131), .QN(n2710)
         );
  DFFR_X1 DR_reg_3_ ( .D(n1152), .CK(i_clk), .RN(n2986), .Q(n3128), .QN(n2709)
         );
  DFFR_X1 DR_reg_2_ ( .D(n1153), .CK(i_clk), .RN(n2986), .Q(n3125), .QN(n2707)
         );
  DFFR_X1 DR_reg_1_ ( .D(n1154), .CK(i_clk), .RN(n2986), .Q(n3122), .QN(n2705)
         );
  DFFR_X1 DR_reg_0_ ( .D(n1155), .CK(i_clk), .RN(n2984), .Q(n3187), .QN(n2703)
         );
  DFFR_X1 DR_reg_31_ ( .D(n1124), .CK(i_clk), .RN(n2999), .Q(n3193), .QN(n2770) );
  DFFR_X1 DR_reg_30_ ( .D(n1125), .CK(i_clk), .RN(n2993), .Q(n3184), .QN(n2736) );
  DFFR_X1 DR_reg_29_ ( .D(n1126), .CK(i_clk), .RN(n2999), .Q(n3182), .QN(n2735) );
  DFFR_X1 DR_reg_28_ ( .D(n1127), .CK(i_clk), .RN(n2998), .Q(n3180), .QN(n2734) );
  DFFR_X1 DR_reg_27_ ( .D(n1128), .CK(i_clk), .RN(n3002), .Q(n3178), .QN(n2733) );
  DFFR_X1 DR_reg_26_ ( .D(n1129), .CK(i_clk), .RN(n2993), .Q(n3176), .QN(n2732) );
  DFFR_X1 DR_reg_25_ ( .D(n1130), .CK(i_clk), .RN(n2999), .Q(n3174), .QN(n2731) );
  DFFR_X1 DR_reg_24_ ( .D(n1131), .CK(i_clk), .RN(n2998), .Q(n3172), .QN(n2730) );
  DFFR_X1 DR_reg_23_ ( .D(n1132), .CK(i_clk), .RN(n2998), .Q(n3170), .QN(n2729) );
  DFFR_X1 DR_reg_22_ ( .D(n1133), .CK(i_clk), .RN(n2995), .Q(n3168), .QN(n2728) );
  DFFR_X1 DR_reg_21_ ( .D(n1134), .CK(i_clk), .RN(n3002), .Q(n3166), .QN(n2727) );
  DFFR_X1 DR_reg_20_ ( .D(n1135), .CK(i_clk), .RN(n2997), .Q(n3164), .QN(n2726) );
  DFFR_X1 DR_reg_19_ ( .D(n1136), .CK(i_clk), .RN(n3004), .Q(n3162), .QN(n2725) );
  DFFR_X1 DR_reg_18_ ( .D(n1137), .CK(i_clk), .RN(n2997), .Q(n3160), .QN(n2724) );
  DFFR_X1 DR_reg_17_ ( .D(n1138), .CK(i_clk), .RN(n2999), .Q(n3158), .QN(n2723) );
  DFFR_X1 DR_reg_16_ ( .D(n1139), .CK(i_clk), .RN(n2996), .Q(n3156), .QN(n2722) );
  DFFR_X1 DR_reg_15_ ( .D(n1140), .CK(i_clk), .RN(n3006), .Q(n3154), .QN(n2721) );
  DFFR_X1 DR_reg_14_ ( .D(n1141), .CK(i_clk), .RN(n2996), .Q(n3152), .QN(n2720) );
  DFFR_X1 DR_reg_13_ ( .D(n1142), .CK(i_clk), .RN(n3008), .Q(n3150), .QN(n2719) );
  DFFR_X1 DR_reg_12_ ( .D(n1143), .CK(i_clk), .RN(n2997), .Q(n3148), .QN(n2718) );
  DFFR_X1 DR_reg_11_ ( .D(n1144), .CK(i_clk), .RN(n2994), .Q(n3146), .QN(n2717) );
  DFFR_X1 DR_reg_10_ ( .D(n1145), .CK(i_clk), .RN(n2997), .Q(n3144), .QN(n2716) );
  DFFR_X1 DR_reg_9_ ( .D(n1146), .CK(i_clk), .RN(n3007), .Q(n3142), .QN(n2715)
         );
  DFFR_X1 DR_reg_8_ ( .D(n1147), .CK(i_clk), .RN(n2996), .Q(n3140), .QN(n2714)
         );
  DFFR_X1 PR_reg_0_ ( .D(n3052), .CK(i_clk), .RN(n2984), .Q(n3053), .QN(n2762)
         );
  DFFR_X1 PR_reg_15_ ( .D(n853), .CK(i_clk), .RN(n3006), .Q(), .QN(n2746) );
  DFFR_X1 PR_reg_13_ ( .D(n855), .CK(i_clk), .RN(n2994), .Q(), .QN(n2744) );
  DFFR_X1 PR_reg_12_ ( .D(n856), .CK(i_clk), .RN(n2995), .Q(), .QN(n2743) );
  DFFR_X1 PR_reg_11_ ( .D(n857), .CK(i_clk), .RN(n3010), .Q(), .QN(n2742) );
  DFFR_X1 PR_reg_16_ ( .D(n852), .CK(i_clk), .RN(n2986), .Q(), .QN(n2747) );
  DFFR_X1 PR_reg_14_ ( .D(n854), .CK(i_clk), .RN(n2986), .Q(), .QN(n2745) );
  DFFR_X1 PR_reg_10_ ( .D(n858), .CK(i_clk), .RN(n2995), .Q(), .QN(n2741) );
  DFFR_X1 PR_reg_26_ ( .D(n842), .CK(i_clk), .RN(n2986), .Q(), .QN(n2757) );
  DFFR_X1 PR_reg_23_ ( .D(n845), .CK(i_clk), .RN(n2986), .Q(), .QN(n2754) );
  DFFR_X1 PR_reg_22_ ( .D(n846), .CK(i_clk), .RN(n2986), .Q(), .QN(n2753) );
  DFFR_X1 PR_reg_30_ ( .D(n838), .CK(i_clk), .RN(n2985), .Q(), .QN(n2761) );
  DFFR_X1 PR_reg_29_ ( .D(n839), .CK(i_clk), .RN(n2985), .Q(), .QN(n2760) );
  DFFR_X1 PR_reg_27_ ( .D(n841), .CK(i_clk), .RN(n2985), .Q(), .QN(n2758) );
  DFFR_X1 PR_reg_25_ ( .D(n843), .CK(i_clk), .RN(n2986), .Q(), .QN(n2756) );
  DFFR_X1 PR_reg_24_ ( .D(n844), .CK(i_clk), .RN(n2986), .Q(), .QN(n2755) );
  DFFR_X1 PR_reg_21_ ( .D(n847), .CK(i_clk), .RN(n3008), .Q(), .QN(n2752) );
  DFFR_X1 PR_reg_20_ ( .D(n848), .CK(i_clk), .RN(n2995), .Q(), .QN(n2751) );
  DFFR_X1 PR_reg_19_ ( .D(n849), .CK(i_clk), .RN(n2995), .Q(), .QN(n2750) );
  DFFR_X1 PR_reg_17_ ( .D(n851), .CK(i_clk), .RN(n3005), .Q(), .QN(n2748) );
  DFFR_X1 PR_reg_18_ ( .D(n850), .CK(i_clk), .RN(n2996), .Q(), .QN(n2749) );
  DFFR_X1 PR_reg_7_ ( .D(n861), .CK(i_clk), .RN(n2995), .Q(), .QN(n2738) );
  DFFR_X1 PR_reg_6_ ( .D(n862), .CK(i_clk), .RN(n2994), .Q(), .QN(n2737) );
  DFFR_X1 PR_reg_8_ ( .D(n860), .CK(i_clk), .RN(n2996), .Q(), .QN(n2739) );
  DFFR_X1 PR_reg_9_ ( .D(n859), .CK(i_clk), .RN(n3007), .Q(), .QN(n2740) );
  DFFR_X1 PR_reg_28_ ( .D(n840), .CK(i_clk), .RN(n2985), .Q(), .QN(n2759) );
  DFFR_X1 PR_reg_1_ ( .D(n3041), .CK(i_clk), .RN(n2985), .Q(n3120), .QN(n2763)
         );
  DFFR_X1 PR_reg_5_ ( .D(n3025), .CK(i_clk), .RN(n3001), .Q(n3132), .QN(n2767)
         );
  DFFR_X1 PR_reg_4_ ( .D(n3026), .CK(i_clk), .RN(n2985), .Q(n3129), .QN(n2766)
         );
  DFFR_X1 PR_reg_3_ ( .D(n3027), .CK(i_clk), .RN(n2985), .Q(n3126), .QN(n2765)
         );
  DFFR_X1 PR_reg_2_ ( .D(n3030), .CK(i_clk), .RN(n2985), .Q(n3123), .QN(n2764)
         );
  DFFR_X1 ct_1_en_1_reg ( .D(n1864), .CK(i_clk), .RN(n3001), .Q(), .QN(n3188)
         );
  DFFR_X1 ready_reg ( .D(n2881), .CK(i_clk), .RN(n3000), .Q(ready), .QN(n3114)
         );
  DFFR_X1 shifted_1_reg_3_ ( .D(n2786), .CK(i_clk), .RN(n3004), .Q(), .QN(
        n3189) );
  DFFR_X1 shifted_1_reg_2_ ( .D(n2785), .CK(i_clk), .RN(n3012), .Q(), .QN(
        n3190) );
  DFFR_X1 shifted_1_reg_1_ ( .D(n2784), .CK(i_clk), .RN(n2987), .Q(), .QN(
        n3191) );
  DFFR_X1 shifted_1_reg_0_ ( .D(n2783), .CK(i_clk), .RN(n3003), .Q(), .QN(
        n3192) );
  DFFR_X1 q_reg_29_ ( .D(n1045), .CK(i_clk), .RN(n2990), .Q(q[29]), .QN(n3225)
         );
  DFFR_X1 q_reg_28_ ( .D(n1046), .CK(i_clk), .RN(n2991), .Q(q[28]), .QN(n3226)
         );
  DFFR_X1 q_reg_27_ ( .D(n1047), .CK(i_clk), .RN(n2989), .Q(q[27]), .QN(n3227)
         );
  DFFR_X1 q_reg_26_ ( .D(n1048), .CK(i_clk), .RN(n2988), .Q(q[26]), .QN(n3228)
         );
  DFFR_X1 q_reg_25_ ( .D(n1049), .CK(i_clk), .RN(n2987), .Q(q[25]), .QN(n3229)
         );
  DFFR_X1 q_reg_24_ ( .D(n1050), .CK(i_clk), .RN(n2987), .Q(q[24]), .QN(n3230)
         );
  DFFR_X1 q_reg_30_ ( .D(n1044), .CK(i_clk), .RN(n2990), .Q(q[30]), .QN(n3224)
         );
  DFFR_X1 nq_reg_30_ ( .D(n1075), .CK(i_clk), .RN(n2990), .Q(nq[30]), .QN(
        n3255) );
  DFFR_X1 nq_reg_29_ ( .D(n1076), .CK(i_clk), .RN(n2990), .Q(nq[29]), .QN(
        n3256) );
  DFFR_X1 nq_reg_28_ ( .D(n1077), .CK(i_clk), .RN(n2991), .Q(nq[28]), .QN(
        n3257) );
  DFFR_X1 nq_reg_27_ ( .D(n1078), .CK(i_clk), .RN(n2989), .Q(nq[27]), .QN(
        n3258) );
  DFFR_X1 nq_reg_26_ ( .D(n1079), .CK(i_clk), .RN(n2988), .Q(nq[26]), .QN(
        n3259) );
  DFFR_X1 nq_reg_25_ ( .D(n1080), .CK(i_clk), .RN(n2987), .Q(nq[25]), .QN(
        n3260) );
  DFFR_X1 nq_reg_24_ ( .D(n1081), .CK(i_clk), .RN(n2987), .Q(nq[24]), .QN(
        n3261) );
  DFFR_X1 q_reg_7_ ( .D(n1067), .CK(i_clk), .RN(n2985), .Q(q[7]), .QN(n3247)
         );
  DFFR_X1 q_reg_6_ ( .D(n1068), .CK(i_clk), .RN(n2990), .Q(q[6]), .QN(n3248)
         );
  DFFR_X1 q_reg_4_ ( .D(n1070), .CK(i_clk), .RN(n2991), .Q(q[4]), .QN(n3250)
         );
  DFFR_X1 q_reg_3_ ( .D(n1071), .CK(i_clk), .RN(n2989), .Q(q[3]), .QN(n3251)
         );
  DFFR_X1 q_reg_2_ ( .D(n1072), .CK(i_clk), .RN(n2989), .Q(q[2]), .QN(n3252)
         );
  DFFR_X1 q_reg_1_ ( .D(n1073), .CK(i_clk), .RN(n2988), .Q(q[1]), .QN(n3253)
         );
  DFFR_X1 q_reg_5_ ( .D(n1069), .CK(i_clk), .RN(n2991), .Q(q[5]), .QN(n3249)
         );
  DFFR_X1 q_reg_11_ ( .D(n1063), .CK(i_clk), .RN(n2989), .Q(q[11]), .QN(n3243)
         );
  DFFR_X1 q_reg_10_ ( .D(n1064), .CK(i_clk), .RN(n2988), .Q(q[10]), .QN(n3244)
         );
  DFFR_X1 q_reg_9_ ( .D(n1065), .CK(i_clk), .RN(n2988), .Q(q[9]), .QN(n3245)
         );
  DFFR_X1 q_reg_8_ ( .D(n1066), .CK(i_clk), .RN(n2984), .Q(q[8]), .QN(n3246)
         );
  DFFR_X1 q_reg_23_ ( .D(n1051), .CK(i_clk), .RN(n2984), .Q(q[23]), .QN(n3231)
         );
  DFFR_X1 q_reg_22_ ( .D(n1052), .CK(i_clk), .RN(n2990), .Q(q[22]), .QN(n3232)
         );
  DFFR_X1 q_reg_21_ ( .D(n1053), .CK(i_clk), .RN(n2990), .Q(q[21]), .QN(n3233)
         );
  DFFR_X1 q_reg_20_ ( .D(n1054), .CK(i_clk), .RN(n2991), .Q(q[20]), .QN(n3234)
         );
  DFFR_X1 q_reg_19_ ( .D(n1055), .CK(i_clk), .RN(n2989), .Q(q[19]), .QN(n3235)
         );
  DFFR_X1 q_reg_18_ ( .D(n1056), .CK(i_clk), .RN(n2988), .Q(q[18]), .QN(n3236)
         );
  DFFR_X1 q_reg_17_ ( .D(n1057), .CK(i_clk), .RN(n2987), .Q(q[17]), .QN(n3237)
         );
  DFFR_X1 q_reg_16_ ( .D(n1058), .CK(i_clk), .RN(n2987), .Q(q[16]), .QN(n3238)
         );
  DFFR_X1 q_reg_15_ ( .D(n1059), .CK(i_clk), .RN(n2984), .Q(q[15]), .QN(n3239)
         );
  DFFR_X1 q_reg_14_ ( .D(n1060), .CK(i_clk), .RN(n2990), .Q(q[14]), .QN(n3240)
         );
  DFFR_X1 q_reg_13_ ( .D(n1061), .CK(i_clk), .RN(n2991), .Q(q[13]), .QN(n3241)
         );
  DFFR_X1 q_reg_12_ ( .D(n1062), .CK(i_clk), .RN(n2991), .Q(q[12]), .QN(n3242)
         );
  DFFR_X1 nq_reg_6_ ( .D(n1099), .CK(i_clk), .RN(n2990), .Q(nq[6]), .QN(n3279)
         );
  DFFR_X1 nq_reg_5_ ( .D(n1100), .CK(i_clk), .RN(n2991), .Q(nq[5]), .QN(n3280)
         );
  DFFR_X1 nq_reg_4_ ( .D(n1101), .CK(i_clk), .RN(n2992), .Q(nq[4]), .QN(n3281)
         );
  DFFR_X1 nq_reg_3_ ( .D(n1102), .CK(i_clk), .RN(n2989), .Q(nq[3]), .QN(n3282)
         );
  DFFR_X1 nq_reg_2_ ( .D(n1103), .CK(i_clk), .RN(n2989), .Q(nq[2]), .QN(n3283)
         );
  DFFR_X1 nq_reg_7_ ( .D(n1098), .CK(i_clk), .RN(n3003), .Q(nq[7]), .QN(n3278)
         );
  DFFR_X1 nq_reg_23_ ( .D(n1082), .CK(i_clk), .RN(n2984), .Q(nq[23]), .QN(
        n3262) );
  DFFR_X1 nq_reg_22_ ( .D(n1083), .CK(i_clk), .RN(n2990), .Q(nq[22]), .QN(
        n3263) );
  DFFR_X1 nq_reg_21_ ( .D(n1084), .CK(i_clk), .RN(n2990), .Q(nq[21]), .QN(
        n3264) );
  DFFR_X1 nq_reg_20_ ( .D(n1085), .CK(i_clk), .RN(n2991), .Q(nq[20]), .QN(
        n3265) );
  DFFR_X1 nq_reg_19_ ( .D(n1086), .CK(i_clk), .RN(n2989), .Q(nq[19]), .QN(
        n3266) );
  DFFR_X1 nq_reg_18_ ( .D(n1087), .CK(i_clk), .RN(n2988), .Q(nq[18]), .QN(
        n3267) );
  DFFR_X1 nq_reg_17_ ( .D(n1088), .CK(i_clk), .RN(n2988), .Q(nq[17]), .QN(
        n3268) );
  DFFR_X1 nq_reg_16_ ( .D(n1089), .CK(i_clk), .RN(n2987), .Q(nq[16]), .QN(
        n3269) );
  DFFR_X1 nq_reg_15_ ( .D(n1090), .CK(i_clk), .RN(n2984), .Q(nq[15]), .QN(
        n3270) );
  DFFR_X1 nq_reg_14_ ( .D(n1091), .CK(i_clk), .RN(n2990), .Q(nq[14]), .QN(
        n3271) );
  DFFR_X1 nq_reg_13_ ( .D(n1092), .CK(i_clk), .RN(n2991), .Q(nq[13]), .QN(
        n3272) );
  DFFR_X1 nq_reg_12_ ( .D(n1093), .CK(i_clk), .RN(n2991), .Q(nq[12]), .QN(
        n3273) );
  DFFR_X1 nq_reg_11_ ( .D(n1094), .CK(i_clk), .RN(n2989), .Q(nq[11]), .QN(
        n3274) );
  DFFR_X1 nq_reg_10_ ( .D(n1095), .CK(i_clk), .RN(n2988), .Q(nq[10]), .QN(
        n3275) );
  DFFR_X1 nq_reg_9_ ( .D(n1096), .CK(i_clk), .RN(n2988), .Q(nq[9]), .QN(n3276)
         );
  DFFR_X1 nq_reg_8_ ( .D(n1097), .CK(i_clk), .RN(n3012), .Q(nq[8]), .QN(n3277)
         );
  DFFR_X1 state_reg_5_ ( .D(n1229), .CK(i_clk), .RN(n2999), .Q(state[5]), .QN(
        n3104) );
  DFFR_X1 state_reg_2_ ( .D(n1226), .CK(i_clk), .RN(n3000), .Q(state[2]), .QN(
        n3108) );
  DFFR_X1 state_reg_1_ ( .D(n1228), .CK(i_clk), .RN(n3000), .Q(state[1]), .QN(
        n3107) );
  DFFR_X1 state_reg_4_ ( .D(n1192), .CK(i_clk), .RN(n3000), .Q(state[4]), .QN(
        n3105) );
  DFFR_X1 state_reg_3_ ( .D(n1225), .CK(i_clk), .RN(n2999), .Q(state[3]), .QN(
        n3109) );
  DFFR_X1 shifted_reg_3_ ( .D(n1187), .CK(i_clk), .RN(n3004), .Q(n2777), .QN(
        n3119) );
  DFFR_X1 shifted_reg_2_ ( .D(n1188), .CK(i_clk), .RN(n3012), .Q(n2778), .QN(
        n3118) );
  DFFR_X1 shifted_reg_1_ ( .D(n1189), .CK(i_clk), .RN(n2987), .Q(n2779), .QN(
        n3117) );
  DFFR_X1 reg_b_reg_5_ ( .D(n1287), .CK(i_clk), .RN(n3001), .Q(reg_b[5]), 
        .QN() );
  DFFR_X1 reg_b_reg_4_ ( .D(n1288), .CK(i_clk), .RN(n3010), .Q(reg_b[4]), 
        .QN() );
  DFFR_X1 reg_b_reg_3_ ( .D(n1289), .CK(i_clk), .RN(n3011), .Q(reg_b[3]), 
        .QN() );
  DFFR_X1 reg_b_reg_2_ ( .D(n1290), .CK(i_clk), .RN(n3011), .Q(reg_b[2]), 
        .QN() );
  DFFR_X1 reg_b_reg_1_ ( .D(n1291), .CK(i_clk), .RN(n2998), .Q(reg_b[1]), 
        .QN() );
  DFFR_X1 reg_b_reg_0_ ( .D(n1292), .CK(i_clk), .RN(n3009), .Q(reg_b[0]), 
        .QN() );
  DFFR_X1 shifted_reg_0_ ( .D(n1190), .CK(i_clk), .RN(n3003), .Q(n2780), .QN(
        n3116) );
  DFFR_X1 PR_reg_31_ ( .D(n3028), .CK(i_clk), .RN(n2984), .Q(n1829), .QN(n3185) );
  DFFR_X1 sdata_reg_0_ ( .D(n2874), .CK(i_clk), .RN(n2984), .Q(sdata[0]), .QN(
        n3115) );
  DFFR_X1 sdata_reg_11_ ( .D(n1175), .CK(i_clk), .RN(n3010), .Q(sdata[11]), 
        .QN(n3145) );
  DFFR_X1 sdata_reg_16_ ( .D(n1170), .CK(i_clk), .RN(n3007), .Q(sdata[16]), 
        .QN(n3155) );
  DFFR_X1 sdata_reg_15_ ( .D(n1171), .CK(i_clk), .RN(n3006), .Q(sdata[15]), 
        .QN(n3153) );
  DFFR_X1 sdata_reg_14_ ( .D(n1172), .CK(i_clk), .RN(n3008), .Q(sdata[14]), 
        .QN(n3151) );
  DFFR_X1 sdata_reg_13_ ( .D(n1173), .CK(i_clk), .RN(n3008), .Q(sdata[13]), 
        .QN(n3149) );
  DFFR_X1 sdata_reg_12_ ( .D(n1174), .CK(i_clk), .RN(n3005), .Q(sdata[12]), 
        .QN(n3147) );
  DFFR_X1 sdata_reg_10_ ( .D(n1176), .CK(i_clk), .RN(n3006), .Q(sdata[10]), 
        .QN(n3143) );
  DFFR_X1 sdata_reg_1_ ( .D(n1185), .CK(i_clk), .RN(n2985), .Q(sdata[1]), .QN(
        n3121) );
  DFFR_X1 sdata_reg_27_ ( .D(n1159), .CK(i_clk), .RN(n3002), .Q(sdata[27]), 
        .QN(n3177) );
  DFFR_X1 sdata_reg_26_ ( .D(n1160), .CK(i_clk), .RN(n3012), .Q(sdata[26]), 
        .QN(n3175) );
  DFFR_X1 sdata_reg_25_ ( .D(n1161), .CK(i_clk), .RN(n2999), .Q(sdata[25]), 
        .QN(n3173) );
  DFFR_X1 sdata_reg_24_ ( .D(n1162), .CK(i_clk), .RN(n3003), .Q(sdata[24]), 
        .QN(n3171) );
  DFFR_X1 sdata_reg_23_ ( .D(n1163), .CK(i_clk), .RN(n3004), .Q(sdata[23]), 
        .QN(n3169) );
  DFFR_X1 sdata_reg_22_ ( .D(n1164), .CK(i_clk), .RN(n3009), .Q(sdata[22]), 
        .QN(n3167) );
  DFFR_X1 sdata_reg_21_ ( .D(n1165), .CK(i_clk), .RN(n3001), .Q(sdata[21]), 
        .QN(n3165) );
  DFFR_X1 sdata_reg_20_ ( .D(n1166), .CK(i_clk), .RN(n3005), .Q(sdata[20]), 
        .QN(n3163) );
  DFFR_X1 sdata_reg_19_ ( .D(n1167), .CK(i_clk), .RN(n3004), .Q(sdata[19]), 
        .QN(n3161) );
  DFFR_X1 sdata_reg_17_ ( .D(n1169), .CK(i_clk), .RN(n2998), .Q(sdata[17]), 
        .QN(n3157) );
  DFFR_X1 sdata_reg_18_ ( .D(n1168), .CK(i_clk), .RN(n3006), .Q(sdata[18]), 
        .QN(n3159) );
  DFFR_X1 sdata_reg_29_ ( .D(n1157), .CK(i_clk), .RN(n2999), .Q(sdata[29]), 
        .QN(n3181) );
  DFFR_X1 sdata_reg_5_ ( .D(n1181), .CK(i_clk), .RN(n2992), .Q(sdata[5]), .QN(
        n3133) );
  DFFR_X1 sdata_reg_4_ ( .D(n1182), .CK(i_clk), .RN(n2986), .Q(sdata[4]), .QN(
        n3130) );
  DFFR_X1 sdata_reg_3_ ( .D(n1183), .CK(i_clk), .RN(n2985), .Q(sdata[3]), .QN(
        n3127) );
  DFFR_X1 sdata_reg_6_ ( .D(n1180), .CK(i_clk), .RN(n2994), .Q(sdata[6]), .QN(
        n3135) );
  DFFR_X1 sdata_reg_7_ ( .D(n1179), .CK(i_clk), .RN(n3010), .Q(sdata[7]), .QN(
        n3137) );
  DFFR_X1 sdata_reg_2_ ( .D(n1184), .CK(i_clk), .RN(n2985), .Q(sdata[2]), .QN(
        n3124) );
  DFFR_X1 sdata_reg_8_ ( .D(n1178), .CK(i_clk), .RN(n3007), .Q(sdata[8]), .QN(
        n3139) );
  DFFR_X1 sdata_reg_9_ ( .D(n1177), .CK(i_clk), .RN(n3007), .Q(sdata[9]), .QN(
        n3141) );
  DFFR_X1 o_remainder_reg_1_ ( .D(n1261), .CK(i_clk), .RN(n3001), .Q(
        o_remainder[1]), .QN(n2638) );
  DFFR_X1 o_remainder_reg_0_ ( .D(n1262), .CK(i_clk), .RN(n3009), .Q(
        o_remainder[0]), .QN(n2637) );
  DFFR_X1 o_remainder_reg_2_ ( .D(n1260), .CK(i_clk), .RN(n3011), .Q(
        o_remainder[2]), .QN(n2639) );
  DFFR_X1 o_quotient_reg_2_ ( .D(n1222), .CK(i_clk), .RN(n3012), .Q(
        o_quotient[2]), .QN(n2671) );
  DFFR_X1 o_quotient_reg_1_ ( .D(n1223), .CK(i_clk), .RN(n3000), .Q(
        o_quotient[1]), .QN(n2670) );
  DFFR_X1 o_quotient_reg_0_ ( .D(n1224), .CK(i_clk), .RN(n3009), .Q(
        o_quotient[0]), .QN(n2669) );
  DFFR_X1 o_quotient_reg_3_ ( .D(n1221), .CK(i_clk), .RN(n3011), .Q(
        o_quotient[3]), .QN(n2672) );
  DFFR_X1 o_remainder_reg_3_ ( .D(n1259), .CK(i_clk), .RN(n3011), .Q(
        o_remainder[3]), .QN(n2640) );
  DFFR_X1 ct_reg_1_ ( .D(n3096), .CK(i_clk), .RN(n3003), .Q(ct[1]), .QN(n938)
         );
  DFFR_X1 ct_reg_0_ ( .D(n3097), .CK(i_clk), .RN(n3003), .Q(ct[0]), .QN(n939)
         );
  DFFR_X1 reg_carry_reg ( .D(n1043), .CK(i_clk), .RN(n2984), .Q(reg_carry), 
        .QN(n940) );
  DFFR_X1 ct_reg_2_ ( .D(n3095), .CK(i_clk), .RN(n2987), .Q(ct[2]), .QN(n937)
         );
  DFFR_X1 o_quotient_reg_5_ ( .D(n1219), .CK(i_clk), .RN(n2992), .Q(
        o_quotient[5]), .QN(n2674) );
  DFFR_X1 o_remainder_reg_5_ ( .D(n1257), .CK(i_clk), .RN(n2992), .Q(
        o_remainder[5]), .QN(n2642) );
  DFFR_X1 o_quotient_reg_4_ ( .D(n1220), .CK(i_clk), .RN(n3010), .Q(
        o_quotient[4]), .QN(n2673) );
  DFFR_X1 o_remainder_reg_4_ ( .D(n1258), .CK(i_clk), .RN(n3010), .Q(
        o_remainder[4]), .QN(n2641) );
  DFFR_X1 ct_reg_3_ ( .D(n3093), .CK(i_clk), .RN(n3012), .Q(ct[3]), .QN(n936)
         );
  DFFR_X1 o_quotient_reg_7_ ( .D(n1217), .CK(i_clk), .RN(n3010), .Q(
        o_quotient[7]), .QN(n2676) );
  DFFR_X1 o_remainder_reg_7_ ( .D(n1255), .CK(i_clk), .RN(n3010), .Q(
        o_remainder[7]), .QN(n2644) );
  DFFR_X1 q_reg_0_ ( .D(n1074), .CK(i_clk), .RN(n2987), .Q(q[0]), .QN(n3254)
         );
  DFFR_X1 nq_reg_1_ ( .D(n1104), .CK(i_clk), .RN(n2988), .Q(n2930), .QN(n3284)
         );
  DFFR_X1 nq_reg_0_ ( .D(n1105), .CK(i_clk), .RN(n2987), .Q(n2931), .QN(n3285)
         );
  DFFR_X1 ct_1_reg_5_ ( .D(n1106), .CK(i_clk), .RN(n2992), .Q(ct_1[5]), .QN(
        n944) );
  DFFR_X1 ct_1_reg_4_ ( .D(n1107), .CK(i_clk), .RN(n3011), .Q(ct_1[4]), .QN(
        n945) );
  DFFR_X1 ct_1_reg_3_ ( .D(n1108), .CK(i_clk), .RN(n3011), .Q(ct_1[3]), .QN(
        n946) );
  DFFR_X1 ct_1_reg_2_ ( .D(n1109), .CK(i_clk), .RN(n3012), .Q(ct_1[2]), .QN(
        n947) );
  DFFR_X1 ct_1_reg_1_ ( .D(n1110), .CK(i_clk), .RN(n2998), .Q(ct_1[1]), .QN(
        n948) );
  DFFR_X1 ct_1_reg_0_ ( .D(n1111), .CK(i_clk), .RN(n3009), .Q(ct_1[0]), .QN(
        n949) );
  DFFR_X1 o_quotient_reg_6_ ( .D(n1218), .CK(i_clk), .RN(n2994), .Q(
        o_quotient[6]), .QN(n2675) );
  DFFR_X1 o_remainder_reg_6_ ( .D(n1256), .CK(i_clk), .RN(n2994), .Q(
        o_remainder[6]), .QN(n2643) );
  DFFR_X1 o_quotient_reg_13_ ( .D(n1211), .CK(i_clk), .RN(n3008), .Q(
        o_quotient[13]), .QN(n2682) );
  DFFR_X1 o_quotient_reg_11_ ( .D(n1213), .CK(i_clk), .RN(n2995), .Q(
        o_quotient[11]), .QN(n2680) );
  DFFR_X1 o_quotient_reg_9_ ( .D(n1215), .CK(i_clk), .RN(n2996), .Q(
        o_quotient[9]), .QN(n2678) );
  DFFR_X1 o_remainder_reg_13_ ( .D(n1249), .CK(i_clk), .RN(n3008), .Q(
        o_remainder[13]), .QN(n2650) );
  DFFR_X1 o_remainder_reg_11_ ( .D(n1251), .CK(i_clk), .RN(n2995), .Q(
        o_remainder[11]), .QN(n2648) );
  DFFR_X1 o_remainder_reg_9_ ( .D(n1253), .CK(i_clk), .RN(n2996), .Q(
        o_remainder[9]), .QN(n2646) );
  DFFR_X1 reg_b_reg_31_ ( .D(n978), .CK(i_clk), .RN(n2984), .Q(reg_b[31]), 
        .QN(n829) );
  DFFR_X1 PR_1_reg_18_ ( .D(n992), .CK(i_clk), .RN(n3006), .Q(PR_1[18]), .QN()
         );
  DFFR_X1 PR_1_reg_16_ ( .D(n994), .CK(i_clk), .RN(n3007), .Q(PR_1[16]), .QN()
         );
  DFFR_X1 PR_1_reg_14_ ( .D(n996), .CK(i_clk), .RN(n3004), .Q(PR_1[14]), .QN()
         );
  DFFR_X1 PR_1_reg_13_ ( .D(n997), .CK(i_clk), .RN(n2993), .Q(PR_1[13]), .QN()
         );
  DFFR_X1 PR_1_reg_11_ ( .D(n999), .CK(i_clk), .RN(n3010), .Q(PR_1[11]), .QN()
         );
  DFFR_X1 PR_1_reg_17_ ( .D(n993), .CK(i_clk), .RN(n2992), .Q(PR_1[17]), .QN()
         );
  DFFR_X1 PR_1_reg_15_ ( .D(n995), .CK(i_clk), .RN(n3011), .Q(PR_1[15]), .QN()
         );
  DFFR_X1 PR_1_reg_12_ ( .D(n998), .CK(i_clk), .RN(n3005), .Q(PR_1[12]), .QN()
         );
  DFFR_X1 ct_reg_4_ ( .D(n3092), .CK(i_clk), .RN(n3012), .Q(ct[4]), .QN(n935)
         );
  DFFR_X1 o_quotient_reg_8_ ( .D(n1216), .CK(i_clk), .RN(n3007), .Q(
        o_quotient[8]), .QN(n2677) );
  DFFR_X1 o_remainder_reg_8_ ( .D(n1254), .CK(i_clk), .RN(n3007), .Q(
        o_remainder[8]), .QN(n2645) );
  DFFR_X1 PR_1_reg_31_ ( .D(n979), .CK(i_clk), .RN(n3001), .Q(PR_1[31]), .QN(
        n870) );
  DFFR_X1 PR_1_reg_30_ ( .D(n980), .CK(i_clk), .RN(n2992), .Q(PR_1[30]), .QN()
         );
  DFFR_X1 PR_1_reg_29_ ( .D(n981), .CK(i_clk), .RN(n2992), .Q(PR_1[29]), .QN()
         );
  DFFR_X1 PR_1_reg_28_ ( .D(n982), .CK(i_clk), .RN(n3002), .Q(PR_1[28]), .QN()
         );
  DFFR_X1 PR_1_reg_27_ ( .D(n983), .CK(i_clk), .RN(n2992), .Q(PR_1[27]), .QN()
         );
  DFFR_X1 PR_1_reg_26_ ( .D(n984), .CK(i_clk), .RN(n3011), .Q(PR_1[26]), .QN()
         );
  DFFR_X1 PR_1_reg_25_ ( .D(n985), .CK(i_clk), .RN(n2993), .Q(PR_1[25]), .QN()
         );
  DFFR_X1 PR_1_reg_24_ ( .D(n986), .CK(i_clk), .RN(n3002), .Q(PR_1[24]), .QN()
         );
  DFFR_X1 PR_1_reg_23_ ( .D(n987), .CK(i_clk), .RN(n3004), .Q(PR_1[23]), .QN()
         );
  DFFR_X1 PR_1_reg_22_ ( .D(n988), .CK(i_clk), .RN(n3009), .Q(PR_1[22]), .QN()
         );
  DFFR_X1 PR_1_reg_21_ ( .D(n989), .CK(i_clk), .RN(n3011), .Q(PR_1[21]), .QN()
         );
  DFFR_X1 PR_1_reg_0_ ( .D(n1010), .CK(i_clk), .RN(n3009), .Q(PR_1[0]), .QN()
         );
  DFFR_X1 PR_1_reg_9_ ( .D(n1001), .CK(i_clk), .RN(n3008), .Q(PR_1[9]), .QN()
         );
  DFFR_X1 PR_1_reg_8_ ( .D(n1002), .CK(i_clk), .RN(n3007), .Q(PR_1[8]), .QN()
         );
  DFFR_X1 PR_1_reg_7_ ( .D(n1003), .CK(i_clk), .RN(n3009), .Q(PR_1[7]), .QN()
         );
  DFFR_X1 PR_1_reg_6_ ( .D(n1004), .CK(i_clk), .RN(n3010), .Q(PR_1[6]), .QN()
         );
  DFFR_X1 PR_1_reg_5_ ( .D(n1005), .CK(i_clk), .RN(n3010), .Q(PR_1[5]), .QN()
         );
  DFFR_X1 PR_1_reg_4_ ( .D(n1006), .CK(i_clk), .RN(n3010), .Q(PR_1[4]), .QN()
         );
  DFFR_X1 PR_1_reg_2_ ( .D(n1008), .CK(i_clk), .RN(n3011), .Q(PR_1[2]), .QN()
         );
  DFFR_X1 PR_1_reg_20_ ( .D(n990), .CK(i_clk), .RN(n3005), .Q(PR_1[20]), .QN()
         );
  DFFR_X1 PR_1_reg_19_ ( .D(n991), .CK(i_clk), .RN(n2993), .Q(PR_1[19]), .QN()
         );
  DFFR_X1 PR_1_reg_10_ ( .D(n1000), .CK(i_clk), .RN(n3006), .Q(PR_1[10]), 
        .QN() );
  DFFR_X1 PR_1_reg_3_ ( .D(n1007), .CK(i_clk), .RN(n3011), .Q(PR_1[3]), .QN()
         );
  DFFR_X1 PR_1_reg_1_ ( .D(n1009), .CK(i_clk), .RN(n3009), .Q(PR_1[1]), .QN()
         );
  DFFR_X1 o_quotient_reg_15_ ( .D(n1209), .CK(i_clk), .RN(n2996), .Q(
        o_quotient[15]), .QN(n2684) );
  DFFR_X1 o_remainder_reg_15_ ( .D(n1247), .CK(i_clk), .RN(n2996), .Q(
        o_remainder[15]), .QN(n2652) );
  DFFR_X1 o_quotient_reg_14_ ( .D(n1210), .CK(i_clk), .RN(n3008), .Q(
        o_quotient[14]), .QN(n2683) );
  DFFR_X1 o_quotient_reg_12_ ( .D(n1212), .CK(i_clk), .RN(n3005), .Q(
        o_quotient[12]), .QN(n2681) );
  DFFR_X1 o_quotient_reg_10_ ( .D(n1214), .CK(i_clk), .RN(n3006), .Q(
        o_quotient[10]), .QN(n2679) );
  DFFR_X1 o_remainder_reg_14_ ( .D(n1248), .CK(i_clk), .RN(n3008), .Q(
        o_remainder[14]), .QN(n2651) );
  DFFR_X1 o_remainder_reg_12_ ( .D(n1250), .CK(i_clk), .RN(n3005), .Q(
        o_remainder[12]), .QN(n2649) );
  DFFR_X1 o_remainder_reg_10_ ( .D(n1252), .CK(i_clk), .RN(n3006), .Q(
        o_remainder[10]), .QN(n2647) );
  DFFR_X1 ct_reg_5_ ( .D(n3094), .CK(i_clk), .RN(n3000), .Q(ct[5]), .QN(n934)
         );
  DFFR_X1 reg_b_reg_11_ ( .D(n1281), .CK(i_clk), .RN(n2994), .Q(reg_b[11]), 
        .QN(n713) );
  DFFR_X1 o_quotient_reg_16_ ( .D(n1208), .CK(i_clk), .RN(n3007), .Q(
        o_quotient[16]), .QN(n2685) );
  DFFR_X1 o_remainder_reg_16_ ( .D(n1246), .CK(i_clk), .RN(n3007), .Q(
        o_remainder[16]), .QN(n2653) );
  DFFR_X1 o_quotient_reg_23_ ( .D(n1201), .CK(i_clk), .RN(n3003), .Q(
        o_quotient[23]), .QN(n2692) );
  DFFR_X1 o_quotient_reg_21_ ( .D(n1203), .CK(i_clk), .RN(n3001), .Q(
        o_quotient[21]), .QN(n2690) );
  DFFR_X1 o_quotient_reg_19_ ( .D(n1205), .CK(i_clk), .RN(n3004), .Q(
        o_quotient[19]), .QN(n2688) );
  DFFR_X1 o_quotient_reg_17_ ( .D(n1207), .CK(i_clk), .RN(n3000), .Q(
        o_quotient[17]), .QN(n2686) );
  DFFR_X1 o_remainder_reg_23_ ( .D(n1239), .CK(i_clk), .RN(n3003), .Q(
        o_remainder[23]), .QN(n2660) );
  DFFR_X1 o_remainder_reg_21_ ( .D(n1241), .CK(i_clk), .RN(n3001), .Q(
        o_remainder[21]), .QN(n2658) );
  DFFR_X1 o_remainder_reg_19_ ( .D(n1243), .CK(i_clk), .RN(n3004), .Q(
        o_remainder[19]), .QN(n2656) );
  DFFR_X1 o_remainder_reg_17_ ( .D(n1245), .CK(i_clk), .RN(n3001), .Q(
        o_remainder[17]), .QN(n2654) );
  DFFR_X1 reg_b_reg_9_ ( .D(n1283), .CK(i_clk), .RN(n3008), .Q(reg_b[9]), .QN(
        n711) );
  DFFR_X1 reg_b_reg_8_ ( .D(n1284), .CK(i_clk), .RN(n3007), .Q(reg_b[8]), .QN(
        n710) );
  DFFR_X1 reg_b_reg_7_ ( .D(n1285), .CK(i_clk), .RN(n3009), .Q(reg_b[7]), .QN(
        n709) );
  DFFR_X1 reg_b_reg_6_ ( .D(n1286), .CK(i_clk), .RN(n2994), .Q(reg_b[6]), .QN(
        n708) );
  DFFR_X1 reg_b_reg_10_ ( .D(n1282), .CK(i_clk), .RN(n3006), .Q(reg_b[10]), 
        .QN(n712) );
  DFFR_X1 o_quotient_reg_27_ ( .D(n1197), .CK(i_clk), .RN(n3002), .Q(
        o_quotient[27]), .QN(n2696) );
  DFFR_X1 o_quotient_reg_25_ ( .D(n1199), .CK(i_clk), .RN(n3000), .Q(
        o_quotient[25]), .QN(n2694) );
  DFFR_X1 o_remainder_reg_27_ ( .D(n1235), .CK(i_clk), .RN(n3002), .Q(
        o_remainder[27]), .QN(n2664) );
  DFFR_X1 o_remainder_reg_25_ ( .D(n1237), .CK(i_clk), .RN(n3001), .Q(
        o_remainder[25]), .QN(n2662) );
  DFFR_X1 o_remainder_reg_31_ ( .D(n1231), .CK(i_clk), .RN(n2998), .Q(
        o_remainder[31]), .QN(n2668) );
  DFFR_X1 o_quotient_reg_29_ ( .D(n1195), .CK(i_clk), .RN(n3000), .Q(
        o_quotient[29]), .QN(n2698) );
  DFFR_X1 o_remainder_reg_29_ ( .D(n1233), .CK(i_clk), .RN(n3001), .Q(
        o_remainder[29]), .QN(n2666) );
  DFFR_X1 o_quotient_reg_31_ ( .D(n1193), .CK(i_clk), .RN(n2998), .Q(
        o_quotient[31]), .QN(n2700) );
  DFFR_X1 reg_b_reg_12_ ( .D(n1280), .CK(i_clk), .RN(n3005), .Q(reg_b[12]), 
        .QN(n714) );
  DFFR_X1 reg_a_reg_31_ ( .D(n2892), .CK(i_clk), .RN(n2984), .Q(reg_a[31]), 
        .QN(n1350) );
  DFFR_X1 o_quotient_reg_24_ ( .D(n1200), .CK(i_clk), .RN(n3003), .Q(
        o_quotient[24]), .QN(n2693) );
  DFFR_X1 o_quotient_reg_22_ ( .D(n1202), .CK(i_clk), .RN(n3009), .Q(
        o_quotient[22]), .QN(n2691) );
  DFFR_X1 o_quotient_reg_20_ ( .D(n1204), .CK(i_clk), .RN(n3005), .Q(
        o_quotient[20]), .QN(n2689) );
  DFFR_X1 o_quotient_reg_18_ ( .D(n1206), .CK(i_clk), .RN(n3006), .Q(
        o_quotient[18]), .QN(n2687) );
  DFFR_X1 o_remainder_reg_24_ ( .D(n1238), .CK(i_clk), .RN(n3003), .Q(
        o_remainder[24]), .QN(n2661) );
  DFFR_X1 o_remainder_reg_22_ ( .D(n1240), .CK(i_clk), .RN(n3009), .Q(
        o_remainder[22]), .QN(n2659) );
  DFFR_X1 o_remainder_reg_20_ ( .D(n1242), .CK(i_clk), .RN(n3004), .Q(
        o_remainder[20]), .QN(n2657) );
  DFFR_X1 o_remainder_reg_18_ ( .D(n1244), .CK(i_clk), .RN(n3005), .Q(
        o_remainder[18]), .QN(n2655) );
  DFFR_X1 reg_a_reg_4_ ( .D(n1038), .CK(i_clk), .RN(n2992), .Q(reg_a[4]), .QN(
        n1769) );
  DFFR_X1 reg_a_reg_3_ ( .D(n1039), .CK(i_clk), .RN(n2989), .Q(reg_a[3]), .QN(
        n1770) );
  DFFR_X1 reg_a_reg_2_ ( .D(n1040), .CK(i_clk), .RN(n2989), .Q(reg_a[2]), .QN(
        n1771) );
  DFFR_X1 reg_a_reg_1_ ( .D(n1041), .CK(i_clk), .RN(n2988), .Q(reg_a[1]), .QN(
        n1772) );
  DFFR_X1 reg_a_reg_0_ ( .D(n1042), .CK(i_clk), .RN(n3005), .Q(reg_a[0]), .QN(
        n1773) );
  DFFR_X1 o_quotient_reg_28_ ( .D(n1196), .CK(i_clk), .RN(n3002), .Q(
        o_quotient[28]), .QN(n2697) );
  DFFR_X1 o_quotient_reg_26_ ( .D(n1198), .CK(i_clk), .RN(n3012), .Q(
        o_quotient[26]), .QN(n2695) );
  DFFR_X1 o_remainder_reg_28_ ( .D(n1234), .CK(i_clk), .RN(n3002), .Q(
        o_remainder[28]), .QN(n2665) );
  DFFR_X1 o_remainder_reg_26_ ( .D(n1236), .CK(i_clk), .RN(n3012), .Q(
        o_remainder[26]), .QN(n2663) );
  DFFR_X1 o_quotient_reg_30_ ( .D(n1194), .CK(i_clk), .RN(n3012), .Q(
        o_quotient[30]), .QN(n2699) );
  DFFR_X1 o_remainder_reg_30_ ( .D(n1232), .CK(i_clk), .RN(n3013), .Q(
        o_remainder[30]), .QN(n2667) );
  DFFR_X1 reg_b_reg_13_ ( .D(n1279), .CK(i_clk), .RN(n2994), .Q(reg_b[13]), 
        .QN(n715) );
  DFFR_X1 reg_a_reg_8_ ( .D(n2791), .CK(i_clk), .RN(n2996), .Q(reg_a[8]), .QN(
        n805) );
  DFFR_X1 reg_a_reg_7_ ( .D(n2792), .CK(i_clk), .RN(n3003), .Q(reg_a[7]), .QN(
        n804) );
  DFFR_X1 reg_a_reg_6_ ( .D(n2793), .CK(i_clk), .RN(n2994), .Q(reg_a[6]), .QN(
        n803) );
  DFFR_X1 reg_a_reg_5_ ( .D(n2794), .CK(i_clk), .RN(n2992), .Q(reg_a[5]), .QN(
        n802) );
  DFFR_X1 reg_a_reg_12_ ( .D(n2808), .CK(i_clk), .RN(n2997), .Q(reg_a[12]), 
        .QN(n809) );
  DFFR_X1 reg_a_reg_11_ ( .D(n2800), .CK(i_clk), .RN(n2994), .Q(reg_a[11]), 
        .QN(n808) );
  DFFR_X1 reg_a_reg_10_ ( .D(n2802), .CK(i_clk), .RN(n2997), .Q(reg_a[10]), 
        .QN(n807) );
  DFFR_X1 reg_a_reg_9_ ( .D(n2803), .CK(i_clk), .RN(n2993), .Q(reg_a[9]), .QN(
        n806) );
  DFFR_X1 reg_a_reg_13_ ( .D(n2805), .CK(i_clk), .RN(n3008), .Q(reg_a[13]), 
        .QN(n810) );
  DFFR_X1 reg_b_reg_14_ ( .D(n1278), .CK(i_clk), .RN(n3004), .Q(reg_b[14]), 
        .QN(n716) );
  DFFR_X1 reg_a_reg_14_ ( .D(n2806), .CK(i_clk), .RN(n2996), .Q(reg_a[14]), 
        .QN(n811) );
  DFFR_X1 reg_b_reg_15_ ( .D(n1277), .CK(i_clk), .RN(n2993), .Q(reg_b[15]), 
        .QN(n717) );
  DFFR_X1 reg_a_reg_15_ ( .D(n2795), .CK(i_clk), .RN(n3006), .Q(reg_a[15]), 
        .QN(n812) );
  DFFR_X1 reg_a_reg_16_ ( .D(n2796), .CK(i_clk), .RN(n2997), .Q(reg_a[16]), 
        .QN(n813) );
  DFFR_X1 reg_b_reg_16_ ( .D(n1276), .CK(i_clk), .RN(n2996), .Q(reg_b[16]), 
        .QN(n718) );
  DFFR_X1 reg_a_reg_17_ ( .D(n2807), .CK(i_clk), .RN(n2999), .Q(reg_a[17]), 
        .QN(n814) );
  DFFR_X1 reg_b_reg_17_ ( .D(n1275), .CK(i_clk), .RN(n3005), .Q(reg_b[17]), 
        .QN(n719) );
  DFFR_X1 reg_b_reg_19_ ( .D(n1273), .CK(i_clk), .RN(n2995), .Q(reg_b[19]), 
        .QN(n721) );
  DFFR_X1 reg_a_reg_18_ ( .D(n2896), .CK(i_clk), .RN(n2997), .Q(reg_a[18]), 
        .QN(n815) );
  DFFR_X1 reg_b_reg_18_ ( .D(n1274), .CK(i_clk), .RN(n2997), .Q(reg_b[18]), 
        .QN(n720) );
  DFFR_X1 reg_b_reg_20_ ( .D(n1272), .CK(i_clk), .RN(n2997), .Q(reg_b[20]), 
        .QN(n722) );
  DFFR_X1 reg_a_reg_19_ ( .D(n2904), .CK(i_clk), .RN(n3004), .Q(reg_a[19]), 
        .QN(n816) );
  DFFR_X1 reg_b_reg_21_ ( .D(n1271), .CK(i_clk), .RN(n3008), .Q(reg_b[21]), 
        .QN(n723) );
  DFFR_X1 reg_a_reg_20_ ( .D(n2894), .CK(i_clk), .RN(n2997), .Q(reg_a[20]), 
        .QN(n817) );
  DFFR_X1 reg_b_reg_22_ ( .D(n1270), .CK(i_clk), .RN(n2995), .Q(reg_b[22]), 
        .QN(n724) );
  DFFR_X1 reg_a_reg_21_ ( .D(n2889), .CK(i_clk), .RN(n3002), .Q(reg_a[21]), 
        .QN(n818) );
  DFFR_X1 reg_b_reg_23_ ( .D(n1269), .CK(i_clk), .RN(n2997), .Q(reg_b[23]), 
        .QN(n725) );
  DFFR_X1 reg_a_reg_22_ ( .D(n2906), .CK(i_clk), .RN(n2995), .Q(reg_a[22]), 
        .QN(n819) );
  DFFR_X1 reg_b_reg_24_ ( .D(n1268), .CK(i_clk), .RN(n3003), .Q(reg_b[24]), 
        .QN(n726) );
  DFFR_X1 reg_a_reg_23_ ( .D(n2910), .CK(i_clk), .RN(n2998), .Q(reg_a[23]), 
        .QN(n820) );
  DFFR_X1 reg_b_reg_25_ ( .D(n1267), .CK(i_clk), .RN(n2993), .Q(reg_b[25]), 
        .QN(n727) );
  DFFR_X1 reg_a_reg_24_ ( .D(n2908), .CK(i_clk), .RN(n2998), .Q(reg_a[24]), 
        .QN(n821) );
  DFFR_X1 reg_b_reg_26_ ( .D(n1266), .CK(i_clk), .RN(n3012), .Q(reg_b[26]), 
        .QN(n728) );
  DFFR_X1 reg_a_reg_25_ ( .D(n2901), .CK(i_clk), .RN(n2999), .Q(reg_a[25]), 
        .QN(n822) );
  DFFR_X1 reg_a_reg_26_ ( .D(n2899), .CK(i_clk), .RN(n2993), .Q(reg_a[26]), 
        .QN(n823) );
  DFFR_X1 reg_b_reg_27_ ( .D(n1265), .CK(i_clk), .RN(n2993), .Q(reg_b[27]), 
        .QN(n729) );
  DFFR_X1 reg_a_reg_29_ ( .D(n2898), .CK(i_clk), .RN(n2999), .Q(reg_a[29]), 
        .QN(n826) );
  DFFR_X1 reg_a_reg_30_ ( .D(n1012), .CK(i_clk), .RN(n3013), .Q(reg_a[30]), 
        .QN(n827) );
  DFFR_X1 reg_a_reg_27_ ( .D(n2801), .CK(i_clk), .RN(n3002), .Q(reg_a[27]), 
        .QN(n824) );
  DFFR_X1 reg_b_reg_28_ ( .D(n1264), .CK(i_clk), .RN(n2998), .Q(reg_b[28]), 
        .QN(n730) );
  DFFR_X1 sdata_reg_31_ ( .D(n1296), .CK(i_clk), .RN(n2999), .Q(sdata[31]), 
        .QN(n3058) );
  DFFR_X1 sdata_reg_30_ ( .D(n1156), .CK(i_clk), .RN(n2991), .Q(sdata[30]), 
        .QN(n3183) );
  DFFR_X1 sdata_reg_28_ ( .D(n1158), .CK(i_clk), .RN(n3002), .Q(sdata[28]), 
        .QN(n3179) );
  DFFR_X1 reg_a_reg_28_ ( .D(n1014), .CK(i_clk), .RN(n2998), .Q(reg_a[28]), 
        .QN(n825) );
  DFFR_X1 reg_b_reg_29_ ( .D(n1263), .CK(i_clk), .RN(n2993), .Q(reg_b[29]), 
        .QN(n731) );
  DFFR_X1 reg_b_reg_30_ ( .D(n1297), .CK(i_clk), .RN(n2993), .Q(reg_b[30]), 
        .QN(n701) );
  NOR2_X2 U2114 ( .A1(nqp1[4]), .A2(n2948), .ZN(n2528) );
  BUF_X1 U2115 ( .A(n2941), .Z(n2942) );
  BUF_X1 U2116 ( .A(n2357), .Z(n2966) );
  AOI211_X1 U2117 ( .C1(n3099), .C2(n3113), .A(n2318), .B(n2319), .ZN(n2311)
         );
  OR2_X1 U2118 ( .A1(n2409), .A2(n3110), .ZN(n2787) );
  AND2_X1 U2119 ( .A1(n2319), .A2(n2451), .ZN(n2788) );
  OR2_X1 U2120 ( .A1(n2939), .A2(n2938), .ZN(n2789) );
  OR2_X1 U2121 ( .A1(n2937), .A2(n2936), .ZN(n2790) );
  BUF_X1 U2122 ( .A(n1034), .Z(n2791) );
  BUF_X1 U2123 ( .A(n1035), .Z(n2792) );
  BUF_X1 U2124 ( .A(n1036), .Z(n2793) );
  BUF_X1 U2125 ( .A(n1037), .Z(n2794) );
  BUF_X1 U2126 ( .A(n1027), .Z(n2795) );
  BUF_X1 U2127 ( .A(n1026), .Z(n2796) );
  NAND2_X2 U2128 ( .A1(n2526), .A2(n2527), .ZN(n1038) );
  NAND2_X2 U2129 ( .A1(n2522), .A2(n2523), .ZN(n1039) );
  INV_X2 U2130 ( .A(i_divisor[30]), .ZN(n3319) );
  BUF_X1 U2131 ( .A(i_dividend[30]), .Z(n2797) );
  INV_X1 U2132 ( .A(n3319), .ZN(n2798) );
  INV_X1 U2133 ( .A(n2798), .ZN(n2799) );
  BUF_X1 U2134 ( .A(n1031), .Z(n2800) );
  BUF_X1 U2135 ( .A(n1015), .Z(n2801) );
  BUF_X1 U2136 ( .A(n1032), .Z(n2802) );
  BUF_X1 U2137 ( .A(n1033), .Z(n2803) );
  BUF_X1 U2138 ( .A(i_dividend[31]), .Z(n2804) );
  BUF_X1 U2139 ( .A(n1029), .Z(n2805) );
  BUF_X1 U2140 ( .A(n1028), .Z(n2806) );
  BUF_X1 U2141 ( .A(n1025), .Z(n2807) );
  BUF_X1 U2142 ( .A(n1030), .Z(n2808) );
  CLKBUF_X1 U2143 ( .A(n2797), .Z(n2809) );
  BUF_X1 U2144 ( .A(i_dividend[26]), .Z(n2810) );
  CLKBUF_X1 U2145 ( .A(n2810), .Z(n2811) );
  BUF_X1 U2146 ( .A(i_dividend[27]), .Z(n2812) );
  BUF_X1 U2147 ( .A(i_divisor[27]), .Z(n2813) );
  CLKBUF_X1 U2148 ( .A(n2812), .Z(n2814) );
  BUF_X1 U2149 ( .A(i_dividend[1]), .Z(n2815) );
  BUF_X1 U2150 ( .A(i_dividend[10]), .Z(n2816) );
  BUF_X1 U2151 ( .A(i_divisor[10]), .Z(n2817) );
  BUF_X1 U2152 ( .A(n2432), .Z(n2818) );
  BUF_X1 U2153 ( .A(i_divisor[12]), .Z(n2819) );
  BUF_X1 U2154 ( .A(n2433), .Z(n2820) );
  BUF_X1 U2155 ( .A(i_divisor[13]), .Z(n2821) );
  BUF_X1 U2156 ( .A(n2434), .Z(n2822) );
  BUF_X1 U2157 ( .A(i_divisor[14]), .Z(n2823) );
  BUF_X1 U2158 ( .A(i_dividend[20]), .Z(n2824) );
  BUF_X1 U2159 ( .A(i_dividend[21]), .Z(n2825) );
  CLKBUF_X1 U2160 ( .A(n2825), .Z(n2826) );
  BUF_X1 U2161 ( .A(i_dividend[22]), .Z(n2827) );
  CLKBUF_X1 U2162 ( .A(n2827), .Z(n2828) );
  BUF_X1 U2163 ( .A(i_dividend[23]), .Z(n2829) );
  CLKBUF_X1 U2164 ( .A(n2829), .Z(n2830) );
  BUF_X1 U2165 ( .A(i_dividend[19]), .Z(n2831) );
  BUF_X1 U2166 ( .A(i_dividend[24]), .Z(n2832) );
  CLKBUF_X1 U2167 ( .A(n2832), .Z(n2833) );
  BUF_X1 U2168 ( .A(i_dividend[25]), .Z(n2834) );
  CLKBUF_X1 U2169 ( .A(n2834), .Z(n2835) );
  BUF_X1 U2170 ( .A(i_dividend[5]), .Z(n2836) );
  BUF_X1 U2171 ( .A(i_divisor[5]), .Z(n2837) );
  CLKBUF_X1 U2172 ( .A(n2836), .Z(n2838) );
  BUF_X1 U2173 ( .A(n3320), .Z(n2839) );
  BUF_X1 U2174 ( .A(i_dividend[29]), .Z(n2840) );
  BUF_X1 U2175 ( .A(i_divisor[29]), .Z(n2841) );
  CLKBUF_X1 U2176 ( .A(n2840), .Z(n2842) );
  BUF_X1 U2177 ( .A(i_dividend[18]), .Z(n2843) );
  BUF_X1 U2178 ( .A(i_dividend[17]), .Z(n2844) );
  BUF_X1 U2179 ( .A(i_divisor[17]), .Z(n2845) );
  CLKBUF_X1 U2180 ( .A(n2824), .Z(n2846) );
  CLKBUF_X1 U2181 ( .A(n2831), .Z(n2847) );
  CLKBUF_X1 U2182 ( .A(n2816), .Z(n2848) );
  CLKBUF_X1 U2183 ( .A(n2815), .Z(n2849) );
  BUF_X1 U2184 ( .A(i_dividend[9]), .Z(n2850) );
  BUF_X1 U2185 ( .A(i_divisor[9]), .Z(n2851) );
  CLKBUF_X1 U2186 ( .A(n2850), .Z(n2852) );
  BUF_X1 U2187 ( .A(i_dividend[8]), .Z(n2853) );
  BUF_X1 U2188 ( .A(i_divisor[8]), .Z(n2854) );
  CLKBUF_X1 U2189 ( .A(n2853), .Z(n2855) );
  BUF_X1 U2190 ( .A(i_dividend[2]), .Z(n2856) );
  CLKBUF_X1 U2191 ( .A(n2856), .Z(n2857) );
  BUF_X1 U2192 ( .A(i_dividend[7]), .Z(n2858) );
  BUF_X1 U2193 ( .A(i_divisor[7]), .Z(n2859) );
  CLKBUF_X1 U2194 ( .A(n2858), .Z(n2860) );
  BUF_X1 U2195 ( .A(i_dividend[6]), .Z(n2861) );
  BUF_X1 U2196 ( .A(i_divisor[6]), .Z(n2862) );
  CLKBUF_X1 U2197 ( .A(n2861), .Z(n2863) );
  BUF_X1 U2198 ( .A(i_dividend[3]), .Z(n2864) );
  CLKBUF_X1 U2199 ( .A(i_divisor[3]), .Z(n2865) );
  CLKBUF_X1 U2200 ( .A(n2864), .Z(n2866) );
  BUF_X1 U2201 ( .A(i_dividend[4]), .Z(n2867) );
  CLKBUF_X1 U2202 ( .A(i_divisor[4]), .Z(n2868) );
  CLKBUF_X1 U2203 ( .A(n2867), .Z(n2869) );
  BUF_X1 U2204 ( .A(n2436), .Z(n2870) );
  BUF_X1 U2205 ( .A(i_divisor[16]), .Z(n2871) );
  BUF_X1 U2206 ( .A(n2431), .Z(n2872) );
  BUF_X1 U2207 ( .A(i_divisor[11]), .Z(n2873) );
  BUF_X1 U2208 ( .A(n1186), .Z(n2874) );
  CLKBUF_X1 U2209 ( .A(i_dividend[0]), .Z(n2875) );
  BUF_X1 U2210 ( .A(n2435), .Z(n2876) );
  BUF_X1 U2211 ( .A(i_divisor[15]), .Z(n2877) );
  NAND2_X2 U2212 ( .A1(n2518), .A2(n2519), .ZN(n1040) );
  CLKBUF_X1 U2213 ( .A(i_divisor[2]), .Z(n2878) );
  CLKBUF_X1 U2214 ( .A(i_dividend[14]), .Z(n2879) );
  NAND2_X2 U2215 ( .A1(n2308), .A2(n2958), .ZN(n1230) );
  INV_X1 U2216 ( .A(n1230), .ZN(n2880) );
  INV_X1 U2217 ( .A(n2880), .ZN(n2881) );
  CLKBUF_X1 U2218 ( .A(i_dividend[16]), .Z(n2882) );
  CLKBUF_X1 U2219 ( .A(n2843), .Z(n2883) );
  CLKBUF_X1 U2220 ( .A(i_dividend[12]), .Z(n2884) );
  CLKBUF_X1 U2221 ( .A(i_dividend[15]), .Z(n2885) );
  CLKBUF_X1 U2222 ( .A(i_dividend[13]), .Z(n2886) );
  CLKBUF_X1 U2223 ( .A(i_dividend[11]), .Z(n2887) );
  CLKBUF_X1 U2224 ( .A(n2844), .Z(n2888) );
  BUF_X1 U2225 ( .A(n1021), .Z(n2889) );
  BUF_X1 U2226 ( .A(i_divisor[21]), .Z(n2890) );
  NAND2_X2 U2227 ( .A1(n2506), .A2(n2507), .ZN(n1042) );
  CLKBUF_X1 U2228 ( .A(i_divisor[0]), .Z(n2891) );
  BUF_X1 U2229 ( .A(n1011), .Z(n2892) );
  CLKBUF_X1 U2230 ( .A(i_divisor[31]), .Z(n2893) );
  BUF_X1 U2231 ( .A(n1022), .Z(n2894) );
  BUF_X1 U2232 ( .A(i_divisor[20]), .Z(n2895) );
  BUF_X1 U2233 ( .A(n1024), .Z(n2896) );
  BUF_X1 U2234 ( .A(i_divisor[18]), .Z(n2897) );
  BUF_X1 U2235 ( .A(n1013), .Z(n2898) );
  BUF_X1 U2236 ( .A(n1016), .Z(n2899) );
  BUF_X1 U2237 ( .A(i_divisor[26]), .Z(n2900) );
  BUF_X1 U2238 ( .A(n1017), .Z(n2901) );
  BUF_X1 U2239 ( .A(i_divisor[25]), .Z(n2902) );
  NAND2_X2 U2240 ( .A1(n2514), .A2(n2515), .ZN(n1041) );
  CLKBUF_X1 U2241 ( .A(i_divisor[1]), .Z(n2903) );
  BUF_X1 U2242 ( .A(n1023), .Z(n2904) );
  BUF_X1 U2243 ( .A(i_divisor[19]), .Z(n2905) );
  BUF_X1 U2244 ( .A(n1020), .Z(n2906) );
  BUF_X1 U2245 ( .A(i_divisor[22]), .Z(n2907) );
  BUF_X1 U2246 ( .A(n1018), .Z(n2908) );
  BUF_X1 U2247 ( .A(i_divisor[24]), .Z(n2909) );
  BUF_X1 U2248 ( .A(n1019), .Z(n2910) );
  BUF_X1 U2249 ( .A(i_divisor[23]), .Z(n2911) );
  INV_X1 U2250 ( .A(i_divisor[28]), .ZN(n2912) );
  INV_X1 U2251 ( .A(n2912), .ZN(n2913) );
  BUF_X1 U2252 ( .A(i_dividend[28]), .Z(n2914) );
  CLKBUF_X1 U2253 ( .A(n2914), .Z(n2915) );
  CLKBUF_X1 U2254 ( .A(n2804), .Z(n2916) );
  OAI221_X1 U2255 ( .B1(n3183), .B2(n2964), .C1(n2799), .C2(n2358), .A(n2450), 
        .ZN(n1156) );
  INV_X2 U2256 ( .A(n2926), .ZN(n2964) );
  OAI221_X1 U2257 ( .B1(n3179), .B2(n2964), .C1(n3321), .C2(n2358), .A(n2448), 
        .ZN(n1158) );
  OAI22_X1 U2258 ( .A1(n2945), .A2(nq[28]), .B1(nqp1[28]), .B2(n2510), .ZN(
        n2603) );
  NAND2_X1 U2259 ( .A1(qp1[30]), .A2(n2357), .ZN(n2922) );
  OAI211_X1 U2260 ( .C1(n2942), .C2(n827), .A(n2608), .B(n2607), .ZN(n1012) );
  OAI22_X1 U2261 ( .A1(n2945), .A2(nq[30]), .B1(nqp1[30]), .B2(n2510), .ZN(
        n2609) );
  OR2_X1 U2262 ( .A1(n2760), .A2(n2975), .ZN(n2917) );
  OR2_X1 U2263 ( .A1(n2941), .A2(n731), .ZN(n2918) );
  NAND3_X1 U2264 ( .A1(n2917), .A2(n2918), .A3(n2400), .ZN(n1263) );
  AND2_X1 U2265 ( .A1(n2969), .A2(PR_1[29]), .ZN(n2919) );
  AND2_X1 U2266 ( .A1(q[29]), .A2(n2967), .ZN(n2920) );
  AND2_X1 U2267 ( .A1(qp1[29]), .A2(n2966), .ZN(n2921) );
  NOR3_X1 U2268 ( .A1(n2919), .A2(n2920), .A3(n2921), .ZN(n2400) );
  NAND2_X1 U2269 ( .A1(n2922), .A2(n2923), .ZN(n1297) );
  NOR2_X1 U2270 ( .A1(n2790), .A2(n2924), .ZN(n2923) );
  NAND2_X1 U2271 ( .A1(n2934), .A2(n2935), .ZN(n2924) );
  INV_X1 U2272 ( .A(n2787), .ZN(n2977) );
  BUF_X1 U2273 ( .A(n2356), .Z(n2967) );
  BUF_X1 U2274 ( .A(n3112), .Z(n2941) );
  INV_X1 U2275 ( .A(n2980), .ZN(n2978) );
  INV_X1 U2276 ( .A(n2980), .ZN(n2979) );
  INV_X1 U2277 ( .A(n2402), .ZN(n2958) );
  BUF_X1 U2278 ( .A(n2511), .Z(n2947) );
  INV_X1 U2279 ( .A(n2403), .ZN(n3057) );
  BUF_X1 U2280 ( .A(n2358), .Z(n2965) );
  BUF_X1 U2281 ( .A(n2510), .Z(n2948) );
  BUF_X1 U2282 ( .A(n2508), .Z(n2949) );
  BUF_X1 U2283 ( .A(n2981), .Z(n2982) );
  BUF_X1 U2284 ( .A(n3091), .Z(n2940) );
  NOR2_X1 U2285 ( .A1(n3098), .A2(n3054), .ZN(n2356) );
  INV_X1 U2286 ( .A(n2366), .ZN(n3112) );
  INV_X1 U2287 ( .A(n2402), .ZN(n2959) );
  INV_X1 U2288 ( .A(n2345), .ZN(n2970) );
  INV_X1 U2289 ( .A(n2974), .ZN(n2971) );
  INV_X1 U2290 ( .A(n2345), .ZN(n2972) );
  BUF_X1 U2291 ( .A(n2457), .Z(n2951) );
  INV_X1 U2292 ( .A(n2788), .ZN(n2953) );
  INV_X1 U2293 ( .A(n2788), .ZN(n2954) );
  INV_X1 U2294 ( .A(n2419), .ZN(n3103) );
  BUF_X1 U2295 ( .A(n2787), .Z(n2980) );
  NOR2_X1 U2296 ( .A1(n2345), .A2(n3113), .ZN(n2366) );
  NAND4_X1 U2297 ( .A1(n2953), .A2(n2958), .A3(n2412), .A4(n2952), .ZN(n2403)
         );
  NOR2_X1 U2298 ( .A1(n977), .A2(n2406), .ZN(n2412) );
  INV_X1 U2299 ( .A(n2928), .ZN(n2969) );
  NOR2_X1 U2300 ( .A1(n2401), .A2(n3098), .ZN(n2357) );
  BUF_X1 U2301 ( .A(n2361), .Z(n2963) );
  BUF_X1 U2302 ( .A(n2363), .Z(n2961) );
  NAND2_X1 U2303 ( .A1(n3113), .A2(n2454), .ZN(n2455) );
  BUF_X1 U2304 ( .A(n2362), .Z(n2962) );
  INV_X1 U2305 ( .A(n2320), .ZN(n3100) );
  BUF_X1 U2306 ( .A(n2512), .Z(n2946) );
  NOR2_X1 U2307 ( .A1(n2610), .A2(n2928), .ZN(n2508) );
  BUF_X1 U2308 ( .A(n2322), .Z(n2981) );
  NOR3_X1 U2309 ( .A1(n2406), .A2(n2973), .A3(n2977), .ZN(n2322) );
  NOR2_X1 U2310 ( .A1(n2401), .A2(n2928), .ZN(n2511) );
  AND2_X1 U2311 ( .A1(n2611), .A2(n2610), .ZN(n2925) );
  AND4_X1 U2312 ( .A1(n2952), .A2(n2940), .A3(n3100), .A4(n3102), .ZN(n2926)
         );
  INV_X1 U2313 ( .A(n2611), .ZN(n3098) );
  INV_X1 U2314 ( .A(sum[4]), .ZN(n3206) );
  INV_X1 U2315 ( .A(sum[5]), .ZN(n3214) );
  NAND2_X1 U2316 ( .A1(n3090), .A2(n2964), .ZN(n2358) );
  INV_X1 U2317 ( .A(n2406), .ZN(n3091) );
  INV_X1 U2318 ( .A(n2465), .ZN(n3081) );
  INV_X1 U2319 ( .A(n2466), .ZN(n3080) );
  INV_X1 U2320 ( .A(n2467), .ZN(n3079) );
  INV_X1 U2321 ( .A(n2468), .ZN(n3078) );
  INV_X1 U2322 ( .A(n2469), .ZN(n3077) );
  INV_X1 U2323 ( .A(n2470), .ZN(n3076) );
  INV_X1 U2324 ( .A(n2471), .ZN(n3075) );
  INV_X1 U2325 ( .A(n2472), .ZN(n3074) );
  INV_X1 U2326 ( .A(n2473), .ZN(n3073) );
  INV_X1 U2327 ( .A(n2474), .ZN(n3072) );
  INV_X1 U2328 ( .A(n2475), .ZN(n3071) );
  INV_X1 U2329 ( .A(n2476), .ZN(n3070) );
  INV_X1 U2330 ( .A(n2477), .ZN(n3069) );
  INV_X1 U2331 ( .A(n2478), .ZN(n3068) );
  INV_X1 U2332 ( .A(n2479), .ZN(n3067) );
  INV_X1 U2333 ( .A(n2480), .ZN(n3066) );
  INV_X1 U2334 ( .A(sum[6]), .ZN(n3213) );
  INV_X1 U2335 ( .A(sum[8]), .ZN(n3198) );
  INV_X1 U2336 ( .A(sum[10]), .ZN(n3217) );
  INV_X1 U2337 ( .A(sum[12]), .ZN(n3202) );
  INV_X1 U2338 ( .A(sum[14]), .ZN(n3209) );
  INV_X1 U2339 ( .A(sum[16]), .ZN(n3194) );
  INV_X1 U2340 ( .A(sum[18]), .ZN(n3219) );
  INV_X1 U2341 ( .A(sum[20]), .ZN(n3204) );
  INV_X1 U2342 ( .A(sum[22]), .ZN(n3211) );
  INV_X1 U2343 ( .A(sum[24]), .ZN(n3196) );
  INV_X1 U2344 ( .A(sum[26]), .ZN(n3215) );
  INV_X1 U2345 ( .A(sum[28]), .ZN(n3200) );
  INV_X1 U2346 ( .A(sum[30]), .ZN(n3056) );
  INV_X1 U2347 ( .A(sum[7]), .ZN(n3199) );
  INV_X1 U2348 ( .A(sum[9]), .ZN(n3218) );
  INV_X1 U2349 ( .A(sum[11]), .ZN(n3203) );
  INV_X1 U2350 ( .A(sum[13]), .ZN(n3210) );
  INV_X1 U2351 ( .A(sum[15]), .ZN(n3195) );
  INV_X1 U2352 ( .A(sum[17]), .ZN(n3220) );
  INV_X1 U2353 ( .A(sum[19]), .ZN(n3205) );
  INV_X1 U2354 ( .A(sum[21]), .ZN(n3212) );
  INV_X1 U2355 ( .A(sum[23]), .ZN(n3197) );
  INV_X1 U2356 ( .A(sum[25]), .ZN(n3216) );
  INV_X1 U2357 ( .A(sum[27]), .ZN(n3201) );
  INV_X1 U2358 ( .A(sum[29]), .ZN(n3208) );
  INV_X1 U2359 ( .A(n2459), .ZN(n3087) );
  INV_X1 U2360 ( .A(n2460), .ZN(n3086) );
  INV_X1 U2361 ( .A(n2461), .ZN(n3085) );
  INV_X1 U2362 ( .A(n2462), .ZN(n3084) );
  INV_X1 U2363 ( .A(n2463), .ZN(n3083) );
  INV_X1 U2364 ( .A(n2464), .ZN(n3082) );
  OR2_X1 U2365 ( .A1(n2610), .A2(n3098), .ZN(n2510) );
  INV_X1 U2366 ( .A(n2481), .ZN(n3065) );
  INV_X1 U2367 ( .A(n2482), .ZN(n3064) );
  INV_X1 U2368 ( .A(n2483), .ZN(n3063) );
  INV_X1 U2369 ( .A(n2484), .ZN(n3062) );
  INV_X1 U2370 ( .A(n2485), .ZN(n3061) );
  INV_X1 U2371 ( .A(n2486), .ZN(n3060) );
  INV_X1 U2372 ( .A(n2487), .ZN(n3059) );
  INV_X1 U2373 ( .A(sum[31]), .ZN(n3055) );
  OR2_X1 U2374 ( .A1(n2975), .A2(n3186), .ZN(n2927) );
  INV_X1 U2375 ( .A(n2319), .ZN(n3102) );
  INV_X1 U2376 ( .A(n2456), .ZN(n3089) );
  INV_X1 U2377 ( .A(n2458), .ZN(n3088) );
  BUF_X1 U2378 ( .A(n2488), .Z(n2950) );
  NOR2_X1 U2379 ( .A1(n2974), .A2(n2319), .ZN(n2419) );
  NAND2_X1 U2380 ( .A1(n2419), .A2(n2413), .ZN(n2414) );
  BUF_X1 U2381 ( .A(n2402), .Z(n2960) );
  INV_X1 U2382 ( .A(sum[2]), .ZN(n3221) );
  INV_X1 U2383 ( .A(sum[1]), .ZN(n3222) );
  INV_X1 U2384 ( .A(sum[3]), .ZN(n3207) );
  INV_X1 U2385 ( .A(n2401), .ZN(n3054) );
  NAND2_X1 U2386 ( .A1(n3186), .A2(n3099), .ZN(n2457) );
  BUF_X1 U2387 ( .A(n2956), .Z(n2957) );
  BUF_X1 U2388 ( .A(n2788), .Z(n2956) );
  BUF_X1 U2389 ( .A(n2788), .Z(n2955) );
  BUF_X1 U2390 ( .A(n2974), .Z(n2973) );
  BUF_X1 U2391 ( .A(n2345), .Z(n2974) );
  OAI21_X1 U2392 ( .B1(n2317), .B2(n3188), .A(n2958), .ZN(n2454) );
  NOR3_X2 U2393 ( .A1(n2408), .A2(n3110), .A3(ct[5]), .ZN(n2320) );
  BUF_X2 U2394 ( .A(n3104), .Z(n2983) );
  OAI21_X1 U2395 ( .B1(n2489), .B2(n2492), .A(n2413), .ZN(n2459) );
  OAI21_X1 U2396 ( .B1(n2489), .B2(n2493), .A(n2413), .ZN(n2460) );
  OAI21_X1 U2397 ( .B1(n2489), .B2(n2494), .A(n2413), .ZN(n2461) );
  OAI21_X1 U2398 ( .B1(n2489), .B2(n2495), .A(n2952), .ZN(n2462) );
  OAI21_X1 U2399 ( .B1(n2489), .B2(n2496), .A(n2413), .ZN(n2463) );
  OAI21_X1 U2400 ( .B1(n2489), .B2(n2497), .A(n2952), .ZN(n2464) );
  NOR2_X1 U2401 ( .A1(n2407), .A2(n3110), .ZN(n2406) );
  NOR2_X1 U2402 ( .A1(n3110), .A2(n2405), .ZN(n2319) );
  OAI21_X1 U2403 ( .B1(n2490), .B2(n2498), .A(n2952), .ZN(n2465) );
  OAI21_X1 U2404 ( .B1(n2491), .B2(n2498), .A(n2952), .ZN(n2466) );
  OAI21_X1 U2405 ( .B1(n2492), .B2(n2498), .A(n2413), .ZN(n2467) );
  OAI21_X1 U2406 ( .B1(n2493), .B2(n2498), .A(n2413), .ZN(n2468) );
  OAI21_X1 U2407 ( .B1(n2494), .B2(n2498), .A(n2413), .ZN(n2469) );
  OAI21_X1 U2408 ( .B1(n2495), .B2(n2498), .A(n2413), .ZN(n2470) );
  OAI21_X1 U2409 ( .B1(n2496), .B2(n2498), .A(n2413), .ZN(n2471) );
  OAI21_X1 U2410 ( .B1(n2497), .B2(n2498), .A(n2413), .ZN(n2472) );
  OAI21_X1 U2411 ( .B1(n2490), .B2(n2499), .A(n2413), .ZN(n2473) );
  OAI21_X1 U2412 ( .B1(n2491), .B2(n2499), .A(n2413), .ZN(n2474) );
  OAI21_X1 U2413 ( .B1(n2492), .B2(n2499), .A(n2413), .ZN(n2475) );
  OAI21_X1 U2414 ( .B1(n2493), .B2(n2499), .A(n2413), .ZN(n2476) );
  OAI21_X1 U2415 ( .B1(n2494), .B2(n2499), .A(n2413), .ZN(n2477) );
  OAI21_X1 U2416 ( .B1(n2495), .B2(n2499), .A(n2413), .ZN(n2478) );
  OAI21_X1 U2417 ( .B1(n2496), .B2(n2499), .A(n2413), .ZN(n2479) );
  OAI21_X1 U2418 ( .B1(n2497), .B2(n2499), .A(n2952), .ZN(n2480) );
  OAI21_X1 U2419 ( .B1(n2489), .B2(n2490), .A(n2413), .ZN(n2456) );
  OAI21_X1 U2420 ( .B1(n2489), .B2(n2491), .A(n2413), .ZN(n2458) );
  OAI21_X1 U2421 ( .B1(n2490), .B2(n2500), .A(n2413), .ZN(n2481) );
  OAI21_X1 U2422 ( .B1(n2491), .B2(n2500), .A(n2952), .ZN(n2482) );
  OAI21_X1 U2423 ( .B1(n2492), .B2(n2500), .A(n2952), .ZN(n2483) );
  OAI21_X1 U2424 ( .B1(n2493), .B2(n2500), .A(n2952), .ZN(n2484) );
  OAI21_X1 U2425 ( .B1(n2494), .B2(n2500), .A(n2952), .ZN(n2485) );
  OAI21_X1 U2426 ( .B1(n2495), .B2(n2500), .A(n2952), .ZN(n2486) );
  OAI21_X1 U2427 ( .B1(n2496), .B2(n2500), .A(n2413), .ZN(n2487) );
  NOR2_X1 U2428 ( .A1(n2410), .A2(n3110), .ZN(n2402) );
  INV_X1 U2429 ( .A(n2502), .ZN(n3110) );
  NOR2_X1 U2430 ( .A1(n2505), .A2(n2409), .ZN(n2611) );
  NOR2_X1 U2431 ( .A1(n2408), .A2(n2926), .ZN(n2362) );
  INV_X1 U2432 ( .A(n2314), .ZN(n3094) );
  AOI22_X1 U2433 ( .A1(sum_ct[5]), .A2(n2310), .B1(n2311), .B2(ct[5]), .ZN(
        n2314) );
  INV_X1 U2434 ( .A(n2315), .ZN(n3093) );
  AOI22_X1 U2435 ( .A1(sum_ct[3]), .A2(n2310), .B1(n2311), .B2(ct[3]), .ZN(
        n2315) );
  OAI22_X1 U2436 ( .A1(n3109), .A2(n2403), .B1(n3057), .B2(n2408), .ZN(n1225)
         );
  OAI22_X1 U2437 ( .A1(n3106), .A2(n2403), .B1(n3057), .B2(n2410), .ZN(n1191)
         );
  NOR2_X1 U2438 ( .A1(n2407), .A2(n2926), .ZN(n2361) );
  OAI22_X1 U2439 ( .A1(n3107), .A2(n2403), .B1(n3057), .B2(n2405), .ZN(n1228)
         );
  OAI22_X1 U2440 ( .A1(n3105), .A2(n2403), .B1(n3057), .B2(n2409), .ZN(n1192)
         );
  OAI22_X1 U2441 ( .A1(n3108), .A2(n2403), .B1(n3057), .B2(n2407), .ZN(n1226)
         );
  OAI22_X1 U2442 ( .A1(n3104), .A2(n2403), .B1(n3057), .B2(n2404), .ZN(n1229)
         );
  OAI22_X1 U2443 ( .A1(n2459), .A2(n3283), .B1(n3087), .B2(n2951), .ZN(n1103)
         );
  OAI22_X1 U2444 ( .A1(n2460), .A2(n3282), .B1(n3086), .B2(n2457), .ZN(n1102)
         );
  OAI22_X1 U2445 ( .A1(n2461), .A2(n3281), .B1(n3085), .B2(n2457), .ZN(n1101)
         );
  NOR2_X1 U2446 ( .A1(n2405), .A2(n2926), .ZN(n2363) );
  NOR2_X1 U2447 ( .A1(n2501), .A2(n2975), .ZN(n2512) );
  BUF_X1 U2448 ( .A(n2413), .Z(n2952) );
  INV_X1 U2449 ( .A(n2317), .ZN(n3113) );
  INV_X1 U2450 ( .A(n2501), .ZN(n3186) );
  OAI21_X1 U2451 ( .B1(n3116), .B2(n2414), .A(n2415), .ZN(n1190) );
  NAND2_X1 U2452 ( .A1(shifted_o[0]), .A2(n3103), .ZN(n2415) );
  OR2_X1 U2453 ( .A1(n2505), .A2(n2410), .ZN(n2928) );
  INV_X1 U2454 ( .A(n2404), .ZN(n3090) );
  OAI21_X1 U2455 ( .B1(n3119), .B2(n2414), .A(n2418), .ZN(n1187) );
  OAI21_X1 U2456 ( .B1(n3118), .B2(n2414), .A(n2417), .ZN(n1188) );
  NAND2_X1 U2457 ( .A1(shifted_o[2]), .A2(n3103), .ZN(n2417) );
  OAI21_X1 U2458 ( .B1(n3117), .B2(n2414), .A(n2416), .ZN(n1189) );
  NAND2_X1 U2459 ( .A1(shifted_o[1]), .A2(n3103), .ZN(n2416) );
  INV_X1 U2460 ( .A(n2313), .ZN(n3095) );
  AOI22_X1 U2461 ( .A1(sum_ct[2]), .A2(n2310), .B1(n2311), .B2(ct[2]), .ZN(
        n2313) );
  INV_X1 U2462 ( .A(n2316), .ZN(n3092) );
  AOI22_X1 U2463 ( .A1(sum_ct[4]), .A2(n2310), .B1(n2311), .B2(ct[4]), .ZN(
        n2316) );
  OR2_X1 U2464 ( .A1(n2977), .A2(n2318), .ZN(n977) );
  INV_X1 U2465 ( .A(n2505), .ZN(n3111) );
  INV_X1 U2466 ( .A(n2353), .ZN(n3025) );
  AOI22_X1 U2467 ( .A1(n2345), .A2(sdata_o[5]), .B1(n3132), .B2(n2972), .ZN(
        n2353) );
  INV_X1 U2468 ( .A(n2352), .ZN(n3026) );
  AOI22_X1 U2469 ( .A1(n2345), .A2(sdata_o[4]), .B1(n3129), .B2(n2970), .ZN(
        n2352) );
  INV_X1 U2470 ( .A(n2351), .ZN(n3027) );
  AOI22_X1 U2471 ( .A1(n2345), .A2(sdata_o[3]), .B1(n3126), .B2(n2972), .ZN(
        n2351) );
  INV_X1 U2472 ( .A(n2350), .ZN(n3030) );
  AOI22_X1 U2473 ( .A1(n2345), .A2(sdata_o[2]), .B1(n3123), .B2(n2970), .ZN(
        n2350) );
  INV_X1 U2474 ( .A(n2349), .ZN(n3041) );
  AOI22_X1 U2475 ( .A1(n2974), .A2(sdata_o[1]), .B1(n3120), .B2(n2971), .ZN(
        n2349) );
  INV_X1 U2476 ( .A(n2348), .ZN(n3052) );
  AOI22_X1 U2477 ( .A1(n2974), .A2(sdata_o[0]), .B1(n3053), .B2(n2971), .ZN(
        n2348) );
  AOI21_X1 U2478 ( .B1(n3102), .B2(n2317), .A(n2311), .ZN(n2310) );
  OAI22_X1 U2479 ( .A1(n2941), .A2(n3188), .B1(n2972), .B2(n2347), .ZN(n1864)
         );
  OAI22_X1 U2480 ( .A1(n2320), .A2(n3192), .B1(n3100), .B2(n3116), .ZN(n2783)
         );
  OAI22_X1 U2481 ( .A1(n2320), .A2(n3191), .B1(n3100), .B2(n3117), .ZN(n2784)
         );
  OAI22_X1 U2482 ( .A1(n2320), .A2(n3190), .B1(n3100), .B2(n3118), .ZN(n2785)
         );
  OAI22_X1 U2483 ( .A1(n2320), .A2(n3189), .B1(n3100), .B2(n3119), .ZN(n2786)
         );
  INV_X1 U2484 ( .A(n2408), .ZN(n3099) );
  NAND2_X1 U2485 ( .A1(n3099), .A2(n2501), .ZN(n2488) );
  INV_X1 U2486 ( .A(sum[0]), .ZN(n3223) );
  INV_X1 U2487 ( .A(n2309), .ZN(n3097) );
  AOI22_X1 U2488 ( .A1(sum_ct[0]), .A2(n2310), .B1(n2311), .B2(ct[0]), .ZN(
        n2309) );
  INV_X1 U2489 ( .A(n2312), .ZN(n3096) );
  AOI22_X1 U2490 ( .A1(sum_ct[1]), .A2(n2310), .B1(n2311), .B2(ct[1]), .ZN(
        n2312) );
  BUF_X1 U2491 ( .A(n3019), .Z(n3016) );
  BUF_X1 U2492 ( .A(n3019), .Z(n3017) );
  BUF_X1 U2493 ( .A(n3019), .Z(n3018) );
  BUF_X1 U2494 ( .A(n3020), .Z(n3015) );
  BUF_X1 U2495 ( .A(n3020), .Z(n3014) );
  INV_X1 U2496 ( .A(n2308), .ZN(o_ready) );
  NOR3_X1 U2497 ( .A1(state[1]), .A2(state[5]), .A3(state[0]), .ZN(n2503) );
  NOR3_X1 U2498 ( .A1(state[3]), .A2(state[4]), .A3(state[2]), .ZN(n2452) );
  OAI221_X1 U2499 ( .B1(n2965), .B2(n3318), .C1(n3058), .C2(n2964), .A(n2360), 
        .ZN(n1296) );
  AOI222_X1 U2500 ( .A1(n2963), .A2(n2916), .B1(sum[31]), .B2(n2962), .C1(
        n2961), .C2(sdata_o[31]), .ZN(n2360) );
  OAI221_X1 U2501 ( .B1(n2965), .B2(n3344), .C1(n2964), .C2(n3133), .A(n2425), 
        .ZN(n1181) );
  AOI222_X1 U2502 ( .A1(n2838), .A2(n2361), .B1(sum[5]), .B2(n2962), .C1(n2961), .C2(sdata_o[5]), .ZN(n2425) );
  OAI221_X1 U2503 ( .B1(n2965), .B2(n3343), .C1(n2964), .C2(n3135), .A(n2426), 
        .ZN(n1180) );
  AOI222_X1 U2504 ( .A1(n2863), .A2(n2963), .B1(sum[6]), .B2(n2362), .C1(n2363), .C2(sdata_o[6]), .ZN(n2426) );
  OAI221_X1 U2505 ( .B1(n2358), .B2(n3345), .C1(n2964), .C2(n3130), .A(n2424), 
        .ZN(n1182) );
  AOI222_X1 U2506 ( .A1(n2869), .A2(n2963), .B1(sum[4]), .B2(n2362), .C1(n2363), .C2(sdata_o[4]), .ZN(n2424) );
  OAI221_X1 U2507 ( .B1(n2358), .B2(n3347), .C1(n2964), .C2(n3124), .A(n2422), 
        .ZN(n1184) );
  AOI222_X1 U2508 ( .A1(n2857), .A2(n2963), .B1(sum[2]), .B2(n2362), .C1(n2363), .C2(sdata_o[2]), .ZN(n2422) );
  OAI221_X1 U2509 ( .B1(n2358), .B2(n3346), .C1(n2964), .C2(n3127), .A(n2423), 
        .ZN(n1183) );
  AOI222_X1 U2510 ( .A1(n2866), .A2(n2963), .B1(sum[3]), .B2(n2362), .C1(n2363), .C2(sdata_o[3]), .ZN(n2423) );
  AOI222_X1 U2511 ( .A1(n2963), .A2(n2809), .B1(sum[30]), .B2(n2962), .C1(
        n2961), .C2(sdata_o[30]), .ZN(n2450) );
  OAI221_X1 U2512 ( .B1(n2965), .B2(n2839), .C1(n3181), .C2(n2964), .A(n2449), 
        .ZN(n1157) );
  AOI222_X1 U2513 ( .A1(n2963), .A2(n2842), .B1(sum[29]), .B2(n2962), .C1(
        n2961), .C2(sdata_o[29]), .ZN(n2449) );
  OAI221_X1 U2514 ( .B1(n2358), .B2(n3342), .C1(n2964), .C2(n3137), .A(n2427), 
        .ZN(n1179) );
  AOI222_X1 U2515 ( .A1(n2860), .A2(n2361), .B1(sum[7]), .B2(n2962), .C1(n2961), .C2(sdata_o[7]), .ZN(n2427) );
  OAI221_X1 U2516 ( .B1(n2358), .B2(n3341), .C1(n2964), .C2(n3139), .A(n2428), 
        .ZN(n1178) );
  AOI222_X1 U2517 ( .A1(n2855), .A2(n2361), .B1(sum[8]), .B2(n2962), .C1(n2961), .C2(sdata_o[8]), .ZN(n2428) );
  OAI221_X1 U2518 ( .B1(n2965), .B2(n3327), .C1(n3167), .C2(n2964), .A(n2442), 
        .ZN(n1164) );
  AOI222_X1 U2519 ( .A1(n2963), .A2(n2828), .B1(sum[22]), .B2(n2962), .C1(
        n2961), .C2(sdata_o[22]), .ZN(n2442) );
  OAI221_X1 U2520 ( .B1(n2965), .B2(n3330), .C1(n3161), .C2(n2964), .A(n2439), 
        .ZN(n1167) );
  AOI222_X1 U2521 ( .A1(n2963), .A2(n2847), .B1(sum[19]), .B2(n2962), .C1(
        n2961), .C2(sdata_o[19]), .ZN(n2439) );
  OAI221_X1 U2522 ( .B1(n2358), .B2(n3332), .C1(n3157), .C2(n2964), .A(n2437), 
        .ZN(n1169) );
  AOI222_X1 U2523 ( .A1(n2963), .A2(n2888), .B1(sum[17]), .B2(n2362), .C1(
        n2363), .C2(sdata_o[17]), .ZN(n2437) );
  OAI221_X1 U2524 ( .B1(n2358), .B2(n3338), .C1(n3145), .C2(n2964), .A(n2872), 
        .ZN(n1175) );
  AOI222_X1 U2525 ( .A1(n2963), .A2(n2887), .B1(sum[11]), .B2(n2962), .C1(
        n2961), .C2(sdata_o[11]), .ZN(n2431) );
  OAI221_X1 U2526 ( .B1(n2358), .B2(n3334), .C1(n3153), .C2(n2964), .A(n2876), 
        .ZN(n1171) );
  AOI222_X1 U2527 ( .A1(n2963), .A2(n2885), .B1(sum[15]), .B2(n2362), .C1(
        n2363), .C2(sdata_o[15]), .ZN(n2435) );
  XNOR2_X1 U2528 ( .A(n1829), .B(n3193), .ZN(n2501) );
  NAND4_X1 U2529 ( .A1(state[2]), .A2(n2503), .A3(n3109), .A4(n3105), .ZN(
        n2408) );
  OAI222_X1 U2530 ( .A1(n2975), .A2(n3185), .B1(n870), .B2(n2928), .C1(n3112), 
        .C2(n829), .ZN(n978) );
  OAI211_X1 U2531 ( .C1(n2942), .C2(n824), .A(n2598), .B(n2599), .ZN(n1015) );
  AOI22_X1 U2532 ( .A1(n2512), .A2(n3178), .B1(n2733), .B2(n2944), .ZN(n2598)
         );
  AOI221_X1 U2533 ( .B1(n2508), .B2(n2813), .C1(n2511), .C2(n3322), .A(n2600), 
        .ZN(n2599) );
  NAND4_X1 U2534 ( .A1(state[4]), .A2(n2503), .A3(n3108), .A4(n3109), .ZN(
        n2410) );
  NAND4_X1 U2535 ( .A1(n2452), .A2(state[5]), .A3(n3106), .A4(n3107), .ZN(
        n2405) );
  AOI22_X1 U2536 ( .A1(n2946), .A2(n3180), .B1(n2734), .B2(n2944), .ZN(n2601)
         );
  AOI221_X1 U2537 ( .B1(n2949), .B2(n2913), .C1(n2947), .C2(n3321), .A(n2603), 
        .ZN(n2602) );
  NAND4_X1 U2538 ( .A1(state[3]), .A2(n2503), .A3(n3108), .A4(n3105), .ZN(
        n2409) );
  AOI222_X1 U2539 ( .A1(n2849), .A2(n2963), .B1(sum[1]), .B2(n2362), .C1(n2363), .C2(sdata_o[1]), .ZN(n2421) );
  AOI222_X1 U2540 ( .A1(n2848), .A2(n2361), .B1(sum[10]), .B2(n2962), .C1(
        n2961), .C2(sdata_o[10]), .ZN(n2430) );
  OAI221_X1 U2541 ( .B1(n2745), .B2(n2975), .C1(n2941), .C2(n716), .A(n2385), 
        .ZN(n1278) );
  AOI222_X1 U2542 ( .A1(n2968), .A2(PR_1[14]), .B1(q[14]), .B2(n2967), .C1(
        qp1[14]), .C2(n2966), .ZN(n2385) );
  OAI221_X1 U2543 ( .B1(n2744), .B2(n2975), .C1(n3112), .C2(n715), .A(n2384), 
        .ZN(n1279) );
  AOI222_X1 U2544 ( .A1(n2968), .A2(PR_1[13]), .B1(q[13]), .B2(n2967), .C1(
        qp1[13]), .C2(n2966), .ZN(n2384) );
  OAI221_X1 U2545 ( .B1(n2743), .B2(n2975), .C1(n2941), .C2(n714), .A(n2383), 
        .ZN(n1280) );
  AOI222_X1 U2546 ( .A1(n2968), .A2(PR_1[12]), .B1(q[12]), .B2(n2967), .C1(
        qp1[12]), .C2(n2966), .ZN(n2383) );
  OAI221_X1 U2547 ( .B1(n2742), .B2(n2975), .C1(n3112), .C2(n713), .A(n2382), 
        .ZN(n1281) );
  AOI222_X1 U2548 ( .A1(n2968), .A2(PR_1[11]), .B1(q[11]), .B2(n2967), .C1(
        qp1[11]), .C2(n2966), .ZN(n2382) );
  OAI221_X1 U2549 ( .B1(n2740), .B2(n2975), .C1(n2941), .C2(n711), .A(n2380), 
        .ZN(n1283) );
  AOI222_X1 U2550 ( .A1(n2968), .A2(PR_1[9]), .B1(q[9]), .B2(n2967), .C1(
        qp1[9]), .C2(n2966), .ZN(n2380) );
  OAI221_X1 U2551 ( .B1(n2739), .B2(n2975), .C1(n3112), .C2(n710), .A(n2379), 
        .ZN(n1284) );
  AOI222_X1 U2552 ( .A1(n2968), .A2(PR_1[8]), .B1(q[8]), .B2(n2356), .C1(
        qp1[8]), .C2(n2357), .ZN(n2379) );
  OAI221_X1 U2553 ( .B1(n2738), .B2(n2975), .C1(n3112), .C2(n709), .A(n2378), 
        .ZN(n1285) );
  AOI222_X1 U2554 ( .A1(n2968), .A2(PR_1[7]), .B1(q[7]), .B2(n2967), .C1(
        qp1[7]), .C2(n2357), .ZN(n2378) );
  OAI221_X1 U2555 ( .B1(n2737), .B2(n2975), .C1(n2941), .C2(n708), .A(n2377), 
        .ZN(n1286) );
  AOI222_X1 U2556 ( .A1(n2968), .A2(PR_1[6]), .B1(q[6]), .B2(n2356), .C1(
        qp1[6]), .C2(n2357), .ZN(n2377) );
  NAND4_X1 U2557 ( .A1(state[1]), .A2(n2452), .A3(n3106), .A4(n3104), .ZN(
        n2407) );
  OAI221_X1 U2558 ( .B1(n2358), .B2(n3349), .C1(n2964), .C2(n3115), .A(n2420), 
        .ZN(n1186) );
  AOI222_X1 U2559 ( .A1(n2875), .A2(n2963), .B1(sum[0]), .B2(n2962), .C1(n2961), .C2(sdata_o[0]), .ZN(n2420) );
  OAI221_X1 U2560 ( .B1(n2504), .B2(n2505), .C1(n2941), .C2(n940), .A(n3098), 
        .ZN(n1043) );
  AOI21_X1 U2561 ( .B1(n2501), .B2(n2410), .A(n3054), .ZN(n2504) );
  OAI221_X1 U2562 ( .B1(n2756), .B2(n2344), .C1(n2941), .C2(n727), .A(n2396), 
        .ZN(n1267) );
  AOI222_X1 U2563 ( .A1(n2969), .A2(PR_1[25]), .B1(q[25]), .B2(n2356), .C1(
        qp1[25]), .C2(n2357), .ZN(n2396) );
  OAI221_X1 U2564 ( .B1(n2752), .B2(n2344), .C1(n2941), .C2(n723), .A(n2392), 
        .ZN(n1271) );
  AOI222_X1 U2565 ( .A1(n2969), .A2(PR_1[21]), .B1(q[21]), .B2(n2967), .C1(
        qp1[21]), .C2(n2966), .ZN(n2392) );
  OAI221_X1 U2566 ( .B1(n2748), .B2(n2344), .C1(n3112), .C2(n719), .A(n2388), 
        .ZN(n1275) );
  AOI222_X1 U2567 ( .A1(n2969), .A2(PR_1[17]), .B1(q[17]), .B2(n2967), .C1(
        qp1[17]), .C2(n2966), .ZN(n2388) );
  OAI22_X1 U2568 ( .A1(n2941), .A2(n1773), .B1(n2927), .B2(n3187), .ZN(n2513)
         );
  OAI22_X1 U2569 ( .A1(n2941), .A2(n1769), .B1(n2927), .B2(n3131), .ZN(n2530)
         );
  OAI22_X1 U2570 ( .A1(n2941), .A2(n1770), .B1(n2927), .B2(n3128), .ZN(n2525)
         );
  OAI22_X1 U2571 ( .A1(n2941), .A2(n1771), .B1(n2927), .B2(n3125), .ZN(n2521)
         );
  OAI22_X1 U2572 ( .A1(n2941), .A2(n1772), .B1(n2927), .B2(n3122), .ZN(n2517)
         );
  OAI221_X1 U2573 ( .B1(n2755), .B2(n2344), .C1(n2941), .C2(n726), .A(n2395), 
        .ZN(n1268) );
  AOI222_X1 U2574 ( .A1(n2969), .A2(PR_1[24]), .B1(q[24]), .B2(n2967), .C1(
        qp1[24]), .C2(n2357), .ZN(n2395) );
  OAI221_X1 U2575 ( .B1(n2754), .B2(n2344), .C1(n2941), .C2(n725), .A(n2394), 
        .ZN(n1269) );
  AOI222_X1 U2576 ( .A1(n2969), .A2(PR_1[23]), .B1(q[23]), .B2(n2967), .C1(
        qp1[23]), .C2(n2357), .ZN(n2394) );
  OAI221_X1 U2577 ( .B1(n2753), .B2(n2344), .C1(n3112), .C2(n724), .A(n2393), 
        .ZN(n1270) );
  AOI222_X1 U2578 ( .A1(n2969), .A2(PR_1[22]), .B1(q[22]), .B2(n2967), .C1(
        qp1[22]), .C2(n2966), .ZN(n2393) );
  OAI221_X1 U2579 ( .B1(n2759), .B2(n2975), .C1(n3112), .C2(n730), .A(n2399), 
        .ZN(n1264) );
  AOI222_X1 U2580 ( .A1(n2969), .A2(PR_1[28]), .B1(q[28]), .B2(n2967), .C1(
        qp1[28]), .C2(n2966), .ZN(n2399) );
  OAI221_X1 U2581 ( .B1(n2757), .B2(n2344), .C1(n2941), .C2(n728), .A(n2397), 
        .ZN(n1266) );
  AOI222_X1 U2582 ( .A1(n2969), .A2(PR_1[26]), .B1(q[26]), .B2(n2967), .C1(
        qp1[26]), .C2(n2966), .ZN(n2397) );
  OAI221_X1 U2583 ( .B1(n2751), .B2(n2344), .C1(n3112), .C2(n722), .A(n2391), 
        .ZN(n1272) );
  AOI222_X1 U2584 ( .A1(n2969), .A2(PR_1[20]), .B1(q[20]), .B2(n2967), .C1(
        qp1[20]), .C2(n2966), .ZN(n2391) );
  OAI221_X1 U2585 ( .B1(n2750), .B2(n2344), .C1(n3112), .C2(n721), .A(n2390), 
        .ZN(n1273) );
  AOI222_X1 U2586 ( .A1(n2969), .A2(PR_1[19]), .B1(q[19]), .B2(n2967), .C1(
        qp1[19]), .C2(n2966), .ZN(n2390) );
  OAI221_X1 U2587 ( .B1(n2749), .B2(n2344), .C1(n2941), .C2(n720), .A(n2389), 
        .ZN(n1274) );
  AOI222_X1 U2588 ( .A1(n2969), .A2(PR_1[18]), .B1(q[18]), .B2(n2967), .C1(
        qp1[18]), .C2(n2966), .ZN(n2389) );
  OAI221_X1 U2589 ( .B1(n2747), .B2(n2344), .C1(n3112), .C2(n718), .A(n2387), 
        .ZN(n1276) );
  AOI222_X1 U2590 ( .A1(n2968), .A2(PR_1[16]), .B1(q[16]), .B2(n2967), .C1(
        qp1[16]), .C2(n2966), .ZN(n2387) );
  OAI221_X1 U2591 ( .B1(n2746), .B2(n2344), .C1(n2941), .C2(n717), .A(n2386), 
        .ZN(n1277) );
  AOI222_X1 U2592 ( .A1(n2968), .A2(PR_1[15]), .B1(q[15]), .B2(n2967), .C1(
        qp1[15]), .C2(n2966), .ZN(n2386) );
  OAI221_X1 U2593 ( .B1(n2741), .B2(n2344), .C1(n3112), .C2(n712), .A(n2381), 
        .ZN(n1282) );
  AOI222_X1 U2594 ( .A1(n2968), .A2(PR_1[10]), .B1(q[10]), .B2(n2356), .C1(
        qp1[10]), .C2(n2357), .ZN(n2381) );
  OAI221_X1 U2595 ( .B1(n2758), .B2(n2344), .C1(n3112), .C2(n729), .A(n2398), 
        .ZN(n1265) );
  AOI222_X1 U2596 ( .A1(n2969), .A2(PR_1[27]), .B1(q[27]), .B2(n2967), .C1(
        qp1[27]), .C2(n2966), .ZN(n2398) );
  OAI221_X1 U2597 ( .B1(n2965), .B2(n3329), .C1(n3163), .C2(n2964), .A(n2440), 
        .ZN(n1166) );
  AOI222_X1 U2598 ( .A1(n2963), .A2(n2846), .B1(sum[20]), .B2(n2962), .C1(
        n2961), .C2(sdata_o[20]), .ZN(n2440) );
  AOI222_X1 U2599 ( .A1(n2361), .A2(n2915), .B1(sum[28]), .B2(n2962), .C1(
        n2961), .C2(sdata_o[28]), .ZN(n2448) );
  OAI221_X1 U2600 ( .B1(n2358), .B2(n3331), .C1(n3159), .C2(n2964), .A(n2438), 
        .ZN(n1168) );
  AOI222_X1 U2601 ( .A1(n2963), .A2(n2883), .B1(sum[18]), .B2(n2962), .C1(
        n2363), .C2(sdata_o[18]), .ZN(n2438) );
  OAI221_X1 U2602 ( .B1(n2358), .B2(n3340), .C1(n2964), .C2(n3141), .A(n2429), 
        .ZN(n1177) );
  AOI222_X1 U2603 ( .A1(n2852), .A2(n2361), .B1(sum[9]), .B2(n2962), .C1(n2961), .C2(sdata_o[9]), .ZN(n2429) );
  OAI221_X1 U2604 ( .B1(n2965), .B2(n3323), .C1(n3175), .C2(n2964), .A(n2446), 
        .ZN(n1160) );
  AOI222_X1 U2605 ( .A1(n2361), .A2(n2811), .B1(sum[26]), .B2(n2962), .C1(
        n2961), .C2(sdata_o[26]), .ZN(n2446) );
  OAI221_X1 U2606 ( .B1(n2965), .B2(n3324), .C1(n3173), .C2(n2964), .A(n2445), 
        .ZN(n1161) );
  AOI222_X1 U2607 ( .A1(n2361), .A2(n2835), .B1(sum[25]), .B2(n2962), .C1(
        n2961), .C2(sdata_o[25]), .ZN(n2445) );
  OAI221_X1 U2608 ( .B1(n2965), .B2(n3326), .C1(n3169), .C2(n2964), .A(n2443), 
        .ZN(n1163) );
  AOI222_X1 U2609 ( .A1(n2361), .A2(n2830), .B1(sum[23]), .B2(n2962), .C1(
        n2961), .C2(sdata_o[23]), .ZN(n2443) );
  OAI221_X1 U2610 ( .B1(n2965), .B2(n3325), .C1(n3171), .C2(n2964), .A(n2444), 
        .ZN(n1162) );
  AOI222_X1 U2611 ( .A1(n2361), .A2(n2833), .B1(sum[24]), .B2(n2962), .C1(
        n2961), .C2(sdata_o[24]), .ZN(n2444) );
  OAI221_X1 U2612 ( .B1(n2965), .B2(n3328), .C1(n3165), .C2(n2964), .A(n2441), 
        .ZN(n1165) );
  AOI222_X1 U2613 ( .A1(n2963), .A2(n2826), .B1(sum[21]), .B2(n2962), .C1(
        n2961), .C2(sdata_o[21]), .ZN(n2441) );
  OAI221_X1 U2614 ( .B1(n2358), .B2(n3333), .C1(n3155), .C2(n2964), .A(n2870), 
        .ZN(n1170) );
  AOI222_X1 U2615 ( .A1(n2963), .A2(n2882), .B1(sum[16]), .B2(n2362), .C1(
        n2363), .C2(sdata_o[16]), .ZN(n2436) );
  OAI221_X1 U2616 ( .B1(n2358), .B2(n3336), .C1(n3149), .C2(n2964), .A(n2820), 
        .ZN(n1173) );
  AOI222_X1 U2617 ( .A1(n2963), .A2(n2886), .B1(sum[13]), .B2(n2362), .C1(
        n2363), .C2(sdata_o[13]), .ZN(n2433) );
  OAI221_X1 U2618 ( .B1(n2358), .B2(n3335), .C1(n3151), .C2(n2964), .A(n2822), 
        .ZN(n1172) );
  AOI222_X1 U2619 ( .A1(n2963), .A2(n2879), .B1(sum[14]), .B2(n2362), .C1(
        n2363), .C2(sdata_o[14]), .ZN(n2434) );
  OAI221_X1 U2620 ( .B1(n2965), .B2(n3337), .C1(n3147), .C2(n2964), .A(n2818), 
        .ZN(n1174) );
  AOI222_X1 U2621 ( .A1(n2963), .A2(n2884), .B1(sum[12]), .B2(n2362), .C1(
        n2363), .C2(sdata_o[12]), .ZN(n2432) );
  OAI221_X1 U2622 ( .B1(n2965), .B2(n3322), .C1(n3177), .C2(n2964), .A(n2447), 
        .ZN(n1159) );
  AOI222_X1 U2623 ( .A1(n2361), .A2(n2814), .B1(sum[27]), .B2(n2962), .C1(
        n2961), .C2(sdata_o[27]), .ZN(n2447) );
  OAI221_X1 U2624 ( .B1(n3091), .B2(n3287), .C1(n2972), .C2(n3183), .A(n2342), 
        .ZN(n980) );
  INV_X1 U2625 ( .A(n2809), .ZN(n3287) );
  AOI22_X1 U2626 ( .A1(n2982), .A2(PR_1[30]), .B1(N294), .B2(n2978), .ZN(n2342) );
  OAI221_X1 U2627 ( .B1(n3091), .B2(n3288), .C1(n2972), .C2(n3181), .A(n2341), 
        .ZN(n981) );
  INV_X1 U2628 ( .A(n2842), .ZN(n3288) );
  AOI22_X1 U2629 ( .A1(n2982), .A2(PR_1[29]), .B1(N293), .B2(n2978), .ZN(n2341) );
  OAI221_X1 U2630 ( .B1(n3091), .B2(n3289), .C1(n2971), .C2(n3179), .A(n2340), 
        .ZN(n982) );
  INV_X1 U2631 ( .A(n2915), .ZN(n3289) );
  AOI22_X1 U2632 ( .A1(n2982), .A2(PR_1[28]), .B1(N292), .B2(n2978), .ZN(n2340) );
  OAI221_X1 U2633 ( .B1(n3091), .B2(n3290), .C1(n2971), .C2(n3177), .A(n2339), 
        .ZN(n983) );
  INV_X1 U2634 ( .A(n2814), .ZN(n3290) );
  AOI22_X1 U2635 ( .A1(n2982), .A2(PR_1[27]), .B1(N291), .B2(n2979), .ZN(n2339) );
  OAI221_X1 U2636 ( .B1(n3091), .B2(n3291), .C1(n2971), .C2(n3175), .A(n2338), 
        .ZN(n984) );
  INV_X1 U2637 ( .A(n2811), .ZN(n3291) );
  AOI22_X1 U2638 ( .A1(n2982), .A2(PR_1[26]), .B1(N290), .B2(n2978), .ZN(n2338) );
  OAI221_X1 U2639 ( .B1(n3091), .B2(n3292), .C1(n2971), .C2(n3173), .A(n2337), 
        .ZN(n985) );
  INV_X1 U2640 ( .A(n2835), .ZN(n3292) );
  AOI22_X1 U2641 ( .A1(n2982), .A2(PR_1[25]), .B1(N289), .B2(n2979), .ZN(n2337) );
  OAI221_X1 U2642 ( .B1(n3091), .B2(n3293), .C1(n2971), .C2(n3171), .A(n2336), 
        .ZN(n986) );
  INV_X1 U2643 ( .A(n2833), .ZN(n3293) );
  AOI22_X1 U2644 ( .A1(n2982), .A2(PR_1[24]), .B1(N288), .B2(n2977), .ZN(n2336) );
  OAI221_X1 U2645 ( .B1(n3091), .B2(n3294), .C1(n2971), .C2(n3169), .A(n2335), 
        .ZN(n987) );
  INV_X1 U2646 ( .A(n2830), .ZN(n3294) );
  AOI22_X1 U2647 ( .A1(n2982), .A2(PR_1[23]), .B1(N287), .B2(n2977), .ZN(n2335) );
  OAI221_X1 U2648 ( .B1(n3091), .B2(n3295), .C1(n2971), .C2(n3167), .A(n2334), 
        .ZN(n988) );
  INV_X1 U2649 ( .A(n2828), .ZN(n3295) );
  AOI22_X1 U2650 ( .A1(n2982), .A2(PR_1[22]), .B1(N286), .B2(n2977), .ZN(n2334) );
  OAI221_X1 U2651 ( .B1(n3091), .B2(n3296), .C1(n2971), .C2(n3165), .A(n2333), 
        .ZN(n989) );
  INV_X1 U2652 ( .A(n2826), .ZN(n3296) );
  AOI22_X1 U2653 ( .A1(n2982), .A2(PR_1[21]), .B1(N285), .B2(n2977), .ZN(n2333) );
  OAI221_X1 U2654 ( .B1(n2940), .B2(n3297), .C1(n2970), .C2(n3163), .A(n2332), 
        .ZN(n990) );
  INV_X1 U2655 ( .A(n2846), .ZN(n3297) );
  AOI22_X1 U2656 ( .A1(n2982), .A2(PR_1[20]), .B1(N284), .B2(n2977), .ZN(n2332) );
  OAI221_X1 U2657 ( .B1(n3091), .B2(n3298), .C1(n2970), .C2(n3161), .A(n2331), 
        .ZN(n991) );
  INV_X1 U2658 ( .A(n2847), .ZN(n3298) );
  AOI22_X1 U2659 ( .A1(n2982), .A2(PR_1[19]), .B1(N283), .B2(n2977), .ZN(n2331) );
  OAI221_X1 U2660 ( .B1(n3091), .B2(n3299), .C1(n2971), .C2(n3159), .A(n2330), 
        .ZN(n992) );
  INV_X1 U2661 ( .A(n2883), .ZN(n3299) );
  AOI22_X1 U2662 ( .A1(n2322), .A2(PR_1[18]), .B1(N282), .B2(n2977), .ZN(n2330) );
  OAI221_X1 U2663 ( .B1(n3091), .B2(n3300), .C1(n2970), .C2(n3157), .A(n2329), 
        .ZN(n993) );
  INV_X1 U2664 ( .A(n2888), .ZN(n3300) );
  AOI22_X1 U2665 ( .A1(n2322), .A2(PR_1[17]), .B1(N281), .B2(n2977), .ZN(n2329) );
  OAI221_X1 U2666 ( .B1(n3091), .B2(n3301), .C1(n2971), .C2(n3155), .A(n2328), 
        .ZN(n994) );
  INV_X1 U2667 ( .A(n2882), .ZN(n3301) );
  AOI22_X1 U2668 ( .A1(n2322), .A2(PR_1[16]), .B1(N280), .B2(n2977), .ZN(n2328) );
  OAI221_X1 U2669 ( .B1(n3091), .B2(n3302), .C1(n2970), .C2(n3153), .A(n2327), 
        .ZN(n995) );
  INV_X1 U2670 ( .A(n2885), .ZN(n3302) );
  AOI22_X1 U2671 ( .A1(n2322), .A2(PR_1[15]), .B1(N279), .B2(n2977), .ZN(n2327) );
  OAI221_X1 U2672 ( .B1(n3091), .B2(n3303), .C1(n2971), .C2(n3151), .A(n2326), 
        .ZN(n996) );
  INV_X1 U2673 ( .A(n2879), .ZN(n3303) );
  AOI22_X1 U2674 ( .A1(n2981), .A2(PR_1[14]), .B1(N278), .B2(n2977), .ZN(n2326) );
  OAI221_X1 U2675 ( .B1(n3091), .B2(n3304), .C1(n2971), .C2(n3149), .A(n2325), 
        .ZN(n997) );
  INV_X1 U2676 ( .A(n2886), .ZN(n3304) );
  AOI22_X1 U2677 ( .A1(n2322), .A2(PR_1[13]), .B1(N277), .B2(n2977), .ZN(n2325) );
  OAI221_X1 U2678 ( .B1(n3091), .B2(n3305), .C1(n2970), .C2(n3147), .A(n2324), 
        .ZN(n998) );
  INV_X1 U2679 ( .A(n2884), .ZN(n3305) );
  AOI22_X1 U2680 ( .A1(n2322), .A2(PR_1[12]), .B1(N276), .B2(n2977), .ZN(n2324) );
  OAI221_X1 U2681 ( .B1(n3091), .B2(n3306), .C1(n2971), .C2(n3145), .A(n2321), 
        .ZN(n999) );
  INV_X1 U2682 ( .A(n2887), .ZN(n3306) );
  AOI22_X1 U2683 ( .A1(n2981), .A2(PR_1[11]), .B1(N275), .B2(n2979), .ZN(n2321) );
  OAI221_X1 U2684 ( .B1(n3091), .B2(n3307), .C1(n2970), .C2(n3143), .A(n2636), 
        .ZN(n1000) );
  INV_X1 U2685 ( .A(n2848), .ZN(n3307) );
  AOI22_X1 U2686 ( .A1(n2981), .A2(PR_1[10]), .B1(N274), .B2(n2977), .ZN(n2636) );
  OAI221_X1 U2687 ( .B1(n3091), .B2(n3286), .C1(n2972), .C2(n3058), .A(n2343), 
        .ZN(n979) );
  AOI22_X1 U2688 ( .A1(n2981), .A2(PR_1[31]), .B1(N295), .B2(n2979), .ZN(n2343) );
  OAI22_X1 U2689 ( .A1(nq[24]), .A2(n2945), .B1(nqp1[24]), .B2(n2948), .ZN(
        n2591) );
  OAI22_X1 U2690 ( .A1(nq[27]), .A2(n2945), .B1(nqp1[27]), .B2(n2510), .ZN(
        n2600) );
  OAI22_X1 U2691 ( .A1(nq[26]), .A2(n2945), .B1(nqp1[26]), .B2(n2510), .ZN(
        n2597) );
  OAI22_X1 U2692 ( .A1(nq[25]), .A2(n2945), .B1(nqp1[25]), .B2(n2510), .ZN(
        n2594) );
  OAI22_X1 U2693 ( .A1(nq[23]), .A2(n2945), .B1(nqp1[23]), .B2(n2510), .ZN(
        n2588) );
  OAI22_X1 U2694 ( .A1(nq[22]), .A2(n2945), .B1(nqp1[22]), .B2(n2510), .ZN(
        n2585) );
  OAI22_X1 U2695 ( .A1(nq[21]), .A2(n2945), .B1(nqp1[21]), .B2(n2510), .ZN(
        n2582) );
  OAI22_X1 U2696 ( .A1(nq[20]), .A2(n2945), .B1(nqp1[20]), .B2(n2510), .ZN(
        n2579) );
  OAI22_X1 U2697 ( .A1(nq[19]), .A2(n2945), .B1(nqp1[19]), .B2(n2510), .ZN(
        n2576) );
  OAI22_X1 U2698 ( .A1(nq[18]), .A2(n2945), .B1(nqp1[18]), .B2(n2510), .ZN(
        n2573) );
  OAI22_X1 U2699 ( .A1(nq[17]), .A2(n2945), .B1(nqp1[17]), .B2(n2510), .ZN(
        n2570) );
  AOI22_X1 U2700 ( .A1(n2946), .A2(n3182), .B1(n2735), .B2(n2943), .ZN(n2604)
         );
  XNOR2_X1 U2701 ( .A(n3058), .B(sdata[30]), .ZN(n2451) );
  NAND2_X1 U2702 ( .A1(n2769), .A2(n3112), .ZN(n2505) );
  NAND4_X1 U2703 ( .A1(n3090), .A2(n2502), .A3(i_start), .A4(n3114), .ZN(n2413) );
  NAND4_X1 U2704 ( .A1(state[0]), .A2(n2452), .A3(n3107), .A4(n3104), .ZN(
        n2404) );
  NOR2_X1 U2705 ( .A1(n941), .A2(state_reg_1_0), .ZN(n2345) );
  OAI22_X1 U2706 ( .A1(n2402), .A2(n2641), .B1(n2958), .B2(n3206), .ZN(n1258)
         );
  OAI22_X1 U2707 ( .A1(n2402), .A2(n2642), .B1(n2958), .B2(n3214), .ZN(n1257)
         );
  OAI22_X1 U2708 ( .A1(n2960), .A2(n2643), .B1(n2958), .B2(n3213), .ZN(n1256)
         );
  OAI22_X1 U2709 ( .A1(n2960), .A2(n2644), .B1(n2958), .B2(n3199), .ZN(n1255)
         );
  OAI22_X1 U2710 ( .A1(n2402), .A2(n2645), .B1(n2958), .B2(n3198), .ZN(n1254)
         );
  OAI22_X1 U2711 ( .A1(n2960), .A2(n2667), .B1(n2958), .B2(n3056), .ZN(n1232)
         );
  OAI22_X1 U2712 ( .A1(n2960), .A2(n2646), .B1(n2959), .B2(n3218), .ZN(n1253)
         );
  OAI22_X1 U2713 ( .A1(n2960), .A2(n2647), .B1(n2959), .B2(n3217), .ZN(n1252)
         );
  OAI22_X1 U2714 ( .A1(n2960), .A2(n2648), .B1(n2959), .B2(n3203), .ZN(n1251)
         );
  OAI22_X1 U2715 ( .A1(n2960), .A2(n2649), .B1(n2959), .B2(n3202), .ZN(n1250)
         );
  OAI22_X1 U2716 ( .A1(n2960), .A2(n2650), .B1(n2959), .B2(n3210), .ZN(n1249)
         );
  OAI22_X1 U2717 ( .A1(n2960), .A2(n2651), .B1(n2959), .B2(n3209), .ZN(n1248)
         );
  OAI22_X1 U2718 ( .A1(n2960), .A2(n2652), .B1(n2959), .B2(n3195), .ZN(n1247)
         );
  OAI22_X1 U2719 ( .A1(n2960), .A2(n2653), .B1(n2959), .B2(n3194), .ZN(n1246)
         );
  OAI22_X1 U2720 ( .A1(n2960), .A2(n2654), .B1(n2959), .B2(n3220), .ZN(n1245)
         );
  OAI22_X1 U2721 ( .A1(n2960), .A2(n2655), .B1(n2959), .B2(n3219), .ZN(n1244)
         );
  OAI22_X1 U2722 ( .A1(n2960), .A2(n2656), .B1(n2959), .B2(n3205), .ZN(n1243)
         );
  OAI22_X1 U2723 ( .A1(n2960), .A2(n2657), .B1(n2959), .B2(n3204), .ZN(n1242)
         );
  OAI221_X1 U2724 ( .B1(n2940), .B2(n3308), .C1(n2972), .C2(n3141), .A(n2635), 
        .ZN(n1001) );
  INV_X1 U2725 ( .A(n2852), .ZN(n3308) );
  AOI22_X1 U2726 ( .A1(n2981), .A2(PR_1[9]), .B1(N273), .B2(n2979), .ZN(n2635)
         );
  OAI221_X1 U2727 ( .B1(n2940), .B2(n3309), .C1(n2972), .C2(n3139), .A(n2634), 
        .ZN(n1002) );
  INV_X1 U2728 ( .A(n2855), .ZN(n3309) );
  AOI22_X1 U2729 ( .A1(n2981), .A2(PR_1[8]), .B1(N272), .B2(n2979), .ZN(n2634)
         );
  OAI221_X1 U2730 ( .B1(n2940), .B2(n3310), .C1(n2972), .C2(n3137), .A(n2633), 
        .ZN(n1003) );
  INV_X1 U2731 ( .A(n2860), .ZN(n3310) );
  AOI22_X1 U2732 ( .A1(n2981), .A2(PR_1[7]), .B1(N271), .B2(n2978), .ZN(n2633)
         );
  OAI221_X1 U2733 ( .B1(n2940), .B2(n3311), .C1(n2972), .C2(n3135), .A(n2632), 
        .ZN(n1004) );
  INV_X1 U2734 ( .A(n2863), .ZN(n3311) );
  AOI22_X1 U2735 ( .A1(n2981), .A2(PR_1[6]), .B1(N270), .B2(n2979), .ZN(n2632)
         );
  OAI221_X1 U2736 ( .B1(n2940), .B2(n3312), .C1(n2972), .C2(n3133), .A(n2631), 
        .ZN(n1005) );
  INV_X1 U2737 ( .A(n2838), .ZN(n3312) );
  AOI22_X1 U2738 ( .A1(n2981), .A2(PR_1[5]), .B1(N269), .B2(n2978), .ZN(n2631)
         );
  OAI221_X1 U2739 ( .B1(n2940), .B2(n3313), .C1(n2972), .C2(n3130), .A(n2630), 
        .ZN(n1006) );
  INV_X1 U2740 ( .A(n2869), .ZN(n3313) );
  AOI22_X1 U2741 ( .A1(n2981), .A2(PR_1[4]), .B1(N268), .B2(n2979), .ZN(n2630)
         );
  OAI22_X1 U2742 ( .A1(n949), .A2(n2454), .B1(n3223), .B2(n2455), .ZN(n1111)
         );
  OAI22_X1 U2743 ( .A1(n948), .A2(n2454), .B1(n3222), .B2(n2455), .ZN(n1110)
         );
  OAI22_X1 U2744 ( .A1(n947), .A2(n2454), .B1(n3221), .B2(n2455), .ZN(n1109)
         );
  OAI22_X1 U2745 ( .A1(n946), .A2(n2454), .B1(n3207), .B2(n2455), .ZN(n1108)
         );
  OAI22_X1 U2746 ( .A1(n945), .A2(n2454), .B1(n3206), .B2(n2455), .ZN(n1107)
         );
  OAI22_X1 U2747 ( .A1(n944), .A2(n2454), .B1(n3214), .B2(n2455), .ZN(n1106)
         );
  OAI22_X1 U2748 ( .A1(n3081), .A2(n2950), .B1(n3246), .B2(n2465), .ZN(n1066)
         );
  OAI22_X1 U2749 ( .A1(n3080), .A2(n2950), .B1(n3245), .B2(n2466), .ZN(n1065)
         );
  OAI22_X1 U2750 ( .A1(n3079), .A2(n2950), .B1(n3244), .B2(n2467), .ZN(n1064)
         );
  OAI22_X1 U2751 ( .A1(n3078), .A2(n2950), .B1(n3243), .B2(n2468), .ZN(n1063)
         );
  OAI22_X1 U2752 ( .A1(n3077), .A2(n2950), .B1(n3242), .B2(n2469), .ZN(n1062)
         );
  OAI22_X1 U2753 ( .A1(n3076), .A2(n2950), .B1(n3241), .B2(n2470), .ZN(n1061)
         );
  OAI22_X1 U2754 ( .A1(n3075), .A2(n2950), .B1(n3240), .B2(n2471), .ZN(n1060)
         );
  OAI22_X1 U2755 ( .A1(n3074), .A2(n2950), .B1(n3239), .B2(n2472), .ZN(n1059)
         );
  OAI22_X1 U2756 ( .A1(n3073), .A2(n2950), .B1(n3238), .B2(n2473), .ZN(n1058)
         );
  OAI22_X1 U2757 ( .A1(n3072), .A2(n2950), .B1(n3237), .B2(n2474), .ZN(n1057)
         );
  OAI22_X1 U2758 ( .A1(n3071), .A2(n2950), .B1(n3236), .B2(n2475), .ZN(n1056)
         );
  OAI22_X1 U2759 ( .A1(n3070), .A2(n2950), .B1(n3235), .B2(n2476), .ZN(n1055)
         );
  OAI22_X1 U2760 ( .A1(n3069), .A2(n2488), .B1(n3234), .B2(n2477), .ZN(n1054)
         );
  OAI22_X1 U2761 ( .A1(n3068), .A2(n2488), .B1(n3233), .B2(n2478), .ZN(n1053)
         );
  OAI22_X1 U2762 ( .A1(n3067), .A2(n2488), .B1(n3232), .B2(n2479), .ZN(n1052)
         );
  OAI22_X1 U2763 ( .A1(n3066), .A2(n2488), .B1(n3231), .B2(n2480), .ZN(n1051)
         );
  OAI22_X1 U2764 ( .A1(n3087), .A2(n2488), .B1(n3252), .B2(n2459), .ZN(n1072)
         );
  OAI22_X1 U2765 ( .A1(n3086), .A2(n2488), .B1(n3251), .B2(n2460), .ZN(n1071)
         );
  OAI22_X1 U2766 ( .A1(n3085), .A2(n2488), .B1(n3250), .B2(n2461), .ZN(n1070)
         );
  OAI22_X1 U2767 ( .A1(n3084), .A2(n2950), .B1(n3249), .B2(n2462), .ZN(n1069)
         );
  OAI22_X1 U2768 ( .A1(n3083), .A2(n2488), .B1(n3248), .B2(n2463), .ZN(n1068)
         );
  OAI22_X1 U2769 ( .A1(n3082), .A2(n2950), .B1(n3247), .B2(n2464), .ZN(n1067)
         );
  OAI22_X1 U2770 ( .A1(n2970), .A2(n3021), .B1(n2740), .B2(n2973), .ZN(n859)
         );
  INV_X1 U2771 ( .A(sdata_o[9]), .ZN(n3021) );
  OAI22_X1 U2772 ( .A1(n2971), .A2(n3044), .B1(n2748), .B2(n2974), .ZN(n851)
         );
  INV_X1 U2773 ( .A(sdata_o[17]), .ZN(n3044) );
  OAI22_X1 U2774 ( .A1(n2970), .A2(n3048), .B1(n2744), .B2(n2974), .ZN(n855)
         );
  INV_X1 U2775 ( .A(sdata_o[13]), .ZN(n3048) );
  OAI22_X1 U2776 ( .A1(n2970), .A2(n3035), .B1(n2756), .B2(n2974), .ZN(n843)
         );
  INV_X1 U2777 ( .A(sdata_o[25]), .ZN(n3035) );
  OAI22_X1 U2778 ( .A1(n2972), .A2(n3039), .B1(n2752), .B2(n2974), .ZN(n847)
         );
  INV_X1 U2779 ( .A(sdata_o[21]), .ZN(n3039) );
  OAI22_X1 U2780 ( .A1(n3065), .A2(n2488), .B1(n3230), .B2(n2481), .ZN(n1050)
         );
  OAI22_X1 U2781 ( .A1(n3064), .A2(n2488), .B1(n3229), .B2(n2482), .ZN(n1049)
         );
  OAI22_X1 U2782 ( .A1(n3063), .A2(n2488), .B1(n3228), .B2(n2483), .ZN(n1048)
         );
  OAI22_X1 U2783 ( .A1(n3062), .A2(n2488), .B1(n3227), .B2(n2484), .ZN(n1047)
         );
  OAI22_X1 U2784 ( .A1(n3061), .A2(n2488), .B1(n3226), .B2(n2485), .ZN(n1046)
         );
  OAI22_X1 U2785 ( .A1(n3060), .A2(n2488), .B1(n3225), .B2(n2486), .ZN(n1045)
         );
  OAI22_X1 U2786 ( .A1(n3059), .A2(n2488), .B1(n3224), .B2(n2487), .ZN(n1044)
         );
  OAI22_X1 U2787 ( .A1(n2402), .A2(n2668), .B1(n3055), .B2(n2958), .ZN(n1231)
         );
  OAI22_X1 U2788 ( .A1(n2970), .A2(n3022), .B1(n2739), .B2(n2973), .ZN(n860)
         );
  INV_X1 U2789 ( .A(sdata_o[8]), .ZN(n3022) );
  OAI22_X1 U2790 ( .A1(n2971), .A2(n3040), .B1(n2751), .B2(n2974), .ZN(n848)
         );
  INV_X1 U2791 ( .A(sdata_o[20]), .ZN(n3040) );
  OAI22_X1 U2792 ( .A1(n2970), .A2(n3045), .B1(n2747), .B2(n2974), .ZN(n852)
         );
  INV_X1 U2793 ( .A(sdata_o[16]), .ZN(n3045) );
  OAI22_X1 U2794 ( .A1(n2970), .A2(n3049), .B1(n2743), .B2(n2973), .ZN(n856)
         );
  INV_X1 U2795 ( .A(sdata_o[12]), .ZN(n3049) );
  OAI22_X1 U2796 ( .A1(n2972), .A2(n3036), .B1(n2755), .B2(n2974), .ZN(n844)
         );
  INV_X1 U2797 ( .A(sdata_o[24]), .ZN(n3036) );
  OAI22_X1 U2798 ( .A1(n2971), .A2(n3032), .B1(n2759), .B2(n2974), .ZN(n840)
         );
  INV_X1 U2799 ( .A(sdata_o[28]), .ZN(n3032) );
  XNOR2_X1 U2800 ( .A(n2778), .B(state[5]), .ZN(n_1_net__2_) );
  XNOR2_X1 U2801 ( .A(n2779), .B(state[5]), .ZN(n_1_net__1_) );
  XNOR2_X1 U2802 ( .A(n2777), .B(state[5]), .ZN(n_1_net__3_) );
  XNOR2_X1 U2803 ( .A(n2780), .B(state[5]), .ZN(n_1_net__0_) );
  OAI22_X1 U2804 ( .A1(n2970), .A2(n3023), .B1(n2738), .B2(n2973), .ZN(n861)
         );
  INV_X1 U2805 ( .A(sdata_o[7]), .ZN(n3023) );
  OAI22_X1 U2806 ( .A1(n2970), .A2(n3050), .B1(n2742), .B2(n2973), .ZN(n857)
         );
  INV_X1 U2807 ( .A(sdata_o[11]), .ZN(n3050) );
  OAI22_X1 U2808 ( .A1(n2972), .A2(n3042), .B1(n2750), .B2(n2974), .ZN(n849)
         );
  INV_X1 U2809 ( .A(sdata_o[19]), .ZN(n3042) );
  OAI22_X1 U2810 ( .A1(n2970), .A2(n3037), .B1(n2754), .B2(n2974), .ZN(n845)
         );
  INV_X1 U2811 ( .A(sdata_o[23]), .ZN(n3037) );
  OAI22_X1 U2812 ( .A1(n2970), .A2(n3046), .B1(n2746), .B2(n2974), .ZN(n853)
         );
  INV_X1 U2813 ( .A(sdata_o[15]), .ZN(n3046) );
  OAI22_X1 U2814 ( .A1(n2971), .A2(n3033), .B1(n2758), .B2(n2974), .ZN(n841)
         );
  INV_X1 U2815 ( .A(sdata_o[27]), .ZN(n3033) );
  OAI22_X1 U2816 ( .A1(n3089), .A2(n2488), .B1(n3254), .B2(n2456), .ZN(n1074)
         );
  OAI22_X1 U2817 ( .A1(n3088), .A2(n2488), .B1(n3253), .B2(n2458), .ZN(n1073)
         );
  OAI22_X1 U2818 ( .A1(n2970), .A2(n3043), .B1(n2749), .B2(n2974), .ZN(n850)
         );
  INV_X1 U2819 ( .A(sdata_o[18]), .ZN(n3043) );
  OAI22_X1 U2820 ( .A1(n2970), .A2(n3024), .B1(n2737), .B2(n2974), .ZN(n862)
         );
  INV_X1 U2821 ( .A(sdata_o[6]), .ZN(n3024) );
  OAI22_X1 U2822 ( .A1(n2972), .A2(n3051), .B1(n2741), .B2(n2974), .ZN(n858)
         );
  INV_X1 U2823 ( .A(sdata_o[10]), .ZN(n3051) );
  OAI22_X1 U2824 ( .A1(n2971), .A2(n3047), .B1(n2745), .B2(n2974), .ZN(n854)
         );
  INV_X1 U2825 ( .A(sdata_o[14]), .ZN(n3047) );
  OAI22_X1 U2826 ( .A1(n2971), .A2(n3038), .B1(n2753), .B2(n2974), .ZN(n846)
         );
  INV_X1 U2827 ( .A(sdata_o[22]), .ZN(n3038) );
  OAI22_X1 U2828 ( .A1(n2972), .A2(n3034), .B1(n2757), .B2(n2974), .ZN(n842)
         );
  INV_X1 U2829 ( .A(sdata_o[26]), .ZN(n3034) );
  OAI22_X1 U2830 ( .A1(n2972), .A2(n3031), .B1(n2760), .B2(n2974), .ZN(n839)
         );
  INV_X1 U2831 ( .A(sdata_o[29]), .ZN(n3031) );
  OAI22_X1 U2832 ( .A1(n2462), .A2(n3280), .B1(n3084), .B2(n2457), .ZN(n1100)
         );
  OAI22_X1 U2833 ( .A1(n2463), .A2(n3279), .B1(n3083), .B2(n2457), .ZN(n1099)
         );
  OAI22_X1 U2834 ( .A1(n2970), .A2(n3029), .B1(n2761), .B2(n2974), .ZN(n838)
         );
  INV_X1 U2835 ( .A(sdata_o[30]), .ZN(n3029) );
  OAI22_X1 U2836 ( .A1(n2960), .A2(n2658), .B1(n2959), .B2(n3212), .ZN(n1241)
         );
  OAI22_X1 U2837 ( .A1(n2960), .A2(n2659), .B1(n2959), .B2(n3211), .ZN(n1240)
         );
  OAI22_X1 U2838 ( .A1(n2960), .A2(n2660), .B1(n2959), .B2(n3197), .ZN(n1239)
         );
  OAI22_X1 U2839 ( .A1(n2960), .A2(n2661), .B1(n2959), .B2(n3196), .ZN(n1238)
         );
  OAI22_X1 U2840 ( .A1(n2960), .A2(n2662), .B1(n2959), .B2(n3216), .ZN(n1237)
         );
  OAI22_X1 U2841 ( .A1(n2960), .A2(n2663), .B1(n2959), .B2(n3215), .ZN(n1236)
         );
  OAI22_X1 U2842 ( .A1(n2960), .A2(n2664), .B1(n2959), .B2(n3201), .ZN(n1235)
         );
  OAI22_X1 U2843 ( .A1(n2960), .A2(n2665), .B1(n2959), .B2(n3200), .ZN(n1234)
         );
  OAI22_X1 U2844 ( .A1(n2402), .A2(n2666), .B1(n2959), .B2(n3208), .ZN(n1233)
         );
  OAI22_X1 U2845 ( .A1(n2464), .A2(n3278), .B1(n3082), .B2(n2951), .ZN(n1098)
         );
  OAI22_X1 U2846 ( .A1(n2465), .A2(n3277), .B1(n3081), .B2(n2951), .ZN(n1097)
         );
  OAI22_X1 U2847 ( .A1(n2466), .A2(n3276), .B1(n3080), .B2(n2951), .ZN(n1096)
         );
  OAI22_X1 U2848 ( .A1(n2467), .A2(n3275), .B1(n3079), .B2(n2951), .ZN(n1095)
         );
  OAI22_X1 U2849 ( .A1(n2468), .A2(n3274), .B1(n3078), .B2(n2951), .ZN(n1094)
         );
  OAI22_X1 U2850 ( .A1(n2469), .A2(n3273), .B1(n3077), .B2(n2951), .ZN(n1093)
         );
  OAI22_X1 U2851 ( .A1(n2470), .A2(n3272), .B1(n3076), .B2(n2951), .ZN(n1092)
         );
  OAI22_X1 U2852 ( .A1(n2471), .A2(n3271), .B1(n3075), .B2(n2951), .ZN(n1091)
         );
  OAI22_X1 U2853 ( .A1(n2472), .A2(n3270), .B1(n3074), .B2(n2951), .ZN(n1090)
         );
  OAI22_X1 U2854 ( .A1(n2473), .A2(n3269), .B1(n3073), .B2(n2951), .ZN(n1089)
         );
  OAI22_X1 U2855 ( .A1(n2474), .A2(n3268), .B1(n3072), .B2(n2951), .ZN(n1088)
         );
  OAI22_X1 U2856 ( .A1(n2475), .A2(n3267), .B1(n3071), .B2(n2951), .ZN(n1087)
         );
  OAI22_X1 U2857 ( .A1(n2476), .A2(n3266), .B1(n3070), .B2(n2951), .ZN(n1086)
         );
  OAI22_X1 U2858 ( .A1(n2477), .A2(n3265), .B1(n3069), .B2(n2457), .ZN(n1085)
         );
  OAI22_X1 U2859 ( .A1(n2478), .A2(n3264), .B1(n3068), .B2(n2457), .ZN(n1084)
         );
  OAI22_X1 U2860 ( .A1(n2479), .A2(n3263), .B1(n3067), .B2(n2457), .ZN(n1083)
         );
  OAI22_X1 U2861 ( .A1(n2480), .A2(n3262), .B1(n3066), .B2(n2457), .ZN(n1082)
         );
  OAI22_X1 U2862 ( .A1(n2481), .A2(n3261), .B1(n3065), .B2(n2457), .ZN(n1081)
         );
  OAI22_X1 U2863 ( .A1(n2482), .A2(n3260), .B1(n3064), .B2(n2457), .ZN(n1080)
         );
  OAI22_X1 U2864 ( .A1(n2483), .A2(n3259), .B1(n3063), .B2(n2457), .ZN(n1079)
         );
  OAI22_X1 U2865 ( .A1(n2484), .A2(n3258), .B1(n3062), .B2(n2457), .ZN(n1078)
         );
  OAI22_X1 U2866 ( .A1(n2485), .A2(n3257), .B1(n3061), .B2(n2457), .ZN(n1077)
         );
  OAI22_X1 U2867 ( .A1(n2486), .A2(n3256), .B1(n3060), .B2(n2457), .ZN(n1076)
         );
  OAI22_X1 U2868 ( .A1(n2487), .A2(n3255), .B1(n3059), .B2(n2457), .ZN(n1075)
         );
  OAI22_X1 U2869 ( .A1(n2978), .A2(n2673), .B1(n2787), .B2(n3206), .ZN(n1220)
         );
  OAI22_X1 U2870 ( .A1(n2978), .A2(n2674), .B1(n2787), .B2(n3214), .ZN(n1219)
         );
  OAI22_X1 U2871 ( .A1(n2979), .A2(n2675), .B1(n2787), .B2(n3213), .ZN(n1218)
         );
  OAI22_X1 U2872 ( .A1(n2978), .A2(n2676), .B1(n2787), .B2(n3199), .ZN(n1217)
         );
  OAI22_X1 U2873 ( .A1(n2978), .A2(n2677), .B1(n2787), .B2(n3198), .ZN(n1216)
         );
  OAI22_X1 U2874 ( .A1(n2979), .A2(n2678), .B1(n2787), .B2(n3218), .ZN(n1215)
         );
  OAI22_X1 U2875 ( .A1(n2978), .A2(n2679), .B1(n2787), .B2(n3217), .ZN(n1214)
         );
  OAI22_X1 U2876 ( .A1(n2979), .A2(n2680), .B1(n2787), .B2(n3203), .ZN(n1213)
         );
  OAI22_X1 U2877 ( .A1(n2978), .A2(n2681), .B1(n2787), .B2(n3202), .ZN(n1212)
         );
  OAI22_X1 U2878 ( .A1(n2978), .A2(n2682), .B1(n2980), .B2(n3210), .ZN(n1211)
         );
  OAI22_X1 U2879 ( .A1(n2979), .A2(n2683), .B1(n2787), .B2(n3209), .ZN(n1210)
         );
  OAI22_X1 U2880 ( .A1(n2978), .A2(n2684), .B1(n2980), .B2(n3195), .ZN(n1209)
         );
  OAI22_X1 U2881 ( .A1(n2978), .A2(n2685), .B1(n2787), .B2(n3194), .ZN(n1208)
         );
  OAI22_X1 U2882 ( .A1(n2979), .A2(n2686), .B1(n2980), .B2(n3220), .ZN(n1207)
         );
  OAI22_X1 U2883 ( .A1(n2978), .A2(n2687), .B1(n2787), .B2(n3219), .ZN(n1206)
         );
  OAI22_X1 U2884 ( .A1(n2978), .A2(n2688), .B1(n2980), .B2(n3205), .ZN(n1205)
         );
  OAI22_X1 U2885 ( .A1(n2979), .A2(n2689), .B1(n2787), .B2(n3204), .ZN(n1204)
         );
  OAI22_X1 U2886 ( .A1(n2978), .A2(n2690), .B1(n2980), .B2(n3212), .ZN(n1203)
         );
  OAI22_X1 U2887 ( .A1(n2979), .A2(n2691), .B1(n2787), .B2(n3211), .ZN(n1202)
         );
  OAI22_X1 U2888 ( .A1(n2978), .A2(n2692), .B1(n2980), .B2(n3197), .ZN(n1201)
         );
  OAI22_X1 U2889 ( .A1(n2979), .A2(n2693), .B1(n2980), .B2(n3196), .ZN(n1200)
         );
  OAI22_X1 U2890 ( .A1(n2979), .A2(n2694), .B1(n2980), .B2(n3216), .ZN(n1199)
         );
  OAI22_X1 U2891 ( .A1(n2979), .A2(n2695), .B1(n2787), .B2(n3215), .ZN(n1198)
         );
  OAI22_X1 U2892 ( .A1(n2979), .A2(n2696), .B1(n2787), .B2(n3201), .ZN(n1197)
         );
  OAI22_X1 U2893 ( .A1(n2979), .A2(n2697), .B1(n2787), .B2(n3200), .ZN(n1196)
         );
  OAI22_X1 U2894 ( .A1(n2979), .A2(n2698), .B1(n2787), .B2(n3208), .ZN(n1195)
         );
  OAI22_X1 U2895 ( .A1(n2978), .A2(n2699), .B1(n2787), .B2(n3056), .ZN(n1194)
         );
  OAI22_X1 U2896 ( .A1(n2979), .A2(n2700), .B1(n2787), .B2(n3055), .ZN(n1193)
         );
  OAI221_X1 U2897 ( .B1(n3091), .B2(n3314), .C1(n2972), .C2(n3127), .A(n2629), 
        .ZN(n1007) );
  INV_X1 U2898 ( .A(n2866), .ZN(n3314) );
  AOI22_X1 U2899 ( .A1(n2981), .A2(PR_1[3]), .B1(N267), .B2(n2978), .ZN(n2629)
         );
  OAI221_X1 U2900 ( .B1(n2940), .B2(n3315), .C1(n2972), .C2(n3124), .A(n2628), 
        .ZN(n1008) );
  INV_X1 U2901 ( .A(n2857), .ZN(n3315) );
  AOI22_X1 U2902 ( .A1(n2981), .A2(PR_1[2]), .B1(N266), .B2(n2979), .ZN(n2628)
         );
  OAI221_X1 U2903 ( .B1(n2940), .B2(n3316), .C1(n2972), .C2(n3121), .A(n2627), 
        .ZN(n1009) );
  INV_X1 U2904 ( .A(n2849), .ZN(n3316) );
  AOI22_X1 U2905 ( .A1(n2981), .A2(PR_1[1]), .B1(N265), .B2(n2978), .ZN(n2627)
         );
  OAI221_X1 U2906 ( .B1(n3091), .B2(n3317), .C1(n2972), .C2(n3115), .A(n2626), 
        .ZN(n1010) );
  INV_X1 U2907 ( .A(n2875), .ZN(n3317) );
  AOI22_X1 U2908 ( .A1(n2981), .A2(PR_1[0]), .B1(N264), .B2(n2978), .ZN(n2626)
         );
  NAND2_X1 U2909 ( .A1(state_reg_1_0), .A2(n941), .ZN(n2317) );
  OAI211_X1 U2910 ( .C1(n944), .C2(n2347), .A(n2375), .B(n2376), .ZN(n1287) );
  AOI222_X1 U2911 ( .A1(reg_b[5]), .A2(n2366), .B1(n2969), .B2(PR_1[5]), .C1(
        n2976), .C2(n3132), .ZN(n2376) );
  AOI22_X1 U2912 ( .A1(q[5]), .A2(n2356), .B1(qp1[5]), .B2(n2966), .ZN(n2375)
         );
  OAI211_X1 U2913 ( .C1(n945), .C2(n2347), .A(n2373), .B(n2374), .ZN(n1288) );
  AOI222_X1 U2914 ( .A1(reg_b[4]), .A2(n2366), .B1(n2969), .B2(PR_1[4]), .C1(
        n2976), .C2(n3129), .ZN(n2374) );
  AOI22_X1 U2915 ( .A1(q[4]), .A2(n2356), .B1(qp1[4]), .B2(n2966), .ZN(n2373)
         );
  OAI211_X1 U2916 ( .C1(n946), .C2(n2347), .A(n2371), .B(n2372), .ZN(n1289) );
  AOI222_X1 U2917 ( .A1(reg_b[3]), .A2(n2366), .B1(n2969), .B2(PR_1[3]), .C1(
        n2976), .C2(n3126), .ZN(n2372) );
  AOI22_X1 U2918 ( .A1(q[3]), .A2(n2356), .B1(qp1[3]), .B2(n2966), .ZN(n2371)
         );
  OAI211_X1 U2919 ( .C1(n947), .C2(n2347), .A(n2369), .B(n2370), .ZN(n1290) );
  AOI222_X1 U2920 ( .A1(reg_b[2]), .A2(n2366), .B1(n2969), .B2(PR_1[2]), .C1(
        n2976), .C2(n3123), .ZN(n2370) );
  AOI22_X1 U2921 ( .A1(q[2]), .A2(n2356), .B1(qp1[2]), .B2(n2357), .ZN(n2369)
         );
  OAI211_X1 U2922 ( .C1(n948), .C2(n2347), .A(n2367), .B(n2368), .ZN(n1291) );
  AOI222_X1 U2923 ( .A1(reg_b[1]), .A2(n2366), .B1(n2969), .B2(PR_1[1]), .C1(
        n2976), .C2(n3120), .ZN(n2368) );
  OAI211_X1 U2924 ( .C1(n949), .C2(n2347), .A(n2364), .B(n2365), .ZN(n1292) );
  AOI222_X1 U2925 ( .A1(reg_b[0]), .A2(n2366), .B1(n2969), .B2(PR_1[0]), .C1(
        n2976), .C2(n3053), .ZN(n2365) );
  AOI22_X1 U2926 ( .A1(n2946), .A2(n3184), .B1(n2736), .B2(n2944), .ZN(n2607)
         );
  NAND4_X1 U2927 ( .A1(n2765), .A2(n2766), .A3(n2767), .A4(n3185), .ZN(n2618)
         );
  OAI211_X1 U2928 ( .C1(n2942), .C2(n821), .A(n2589), .B(n2590), .ZN(n1018) );
  AOI22_X1 U2929 ( .A1(n2512), .A2(n3172), .B1(n2730), .B2(n2944), .ZN(n2589)
         );
  AOI221_X1 U2930 ( .B1(n2949), .B2(n2909), .C1(n2947), .C2(n3325), .A(n2591), 
        .ZN(n2590) );
  OAI211_X1 U2931 ( .C1(n2942), .C2(n820), .A(n2586), .B(n2587), .ZN(n1019) );
  AOI22_X1 U2932 ( .A1(n2512), .A2(n3170), .B1(n2729), .B2(n2944), .ZN(n2586)
         );
  AOI221_X1 U2933 ( .B1(n2949), .B2(n2911), .C1(n2947), .C2(n3326), .A(n2588), 
        .ZN(n2587) );
  OAI211_X1 U2934 ( .C1(n2942), .C2(n819), .A(n2583), .B(n2584), .ZN(n1020) );
  AOI22_X1 U2935 ( .A1(n2946), .A2(n3168), .B1(n2728), .B2(n2944), .ZN(n2583)
         );
  AOI221_X1 U2936 ( .B1(n2949), .B2(n2907), .C1(n2947), .C2(n3327), .A(n2585), 
        .ZN(n2584) );
  OAI211_X1 U2937 ( .C1(n3112), .C2(n818), .A(n2580), .B(n2581), .ZN(n1021) );
  AOI22_X1 U2938 ( .A1(n2512), .A2(n3166), .B1(n2727), .B2(n2944), .ZN(n2580)
         );
  AOI221_X1 U2939 ( .B1(n2508), .B2(n2890), .C1(n2947), .C2(n3328), .A(n2582), 
        .ZN(n2581) );
  OAI211_X1 U2940 ( .C1(n2942), .C2(n823), .A(n2595), .B(n2596), .ZN(n1016) );
  AOI22_X1 U2941 ( .A1(n2946), .A2(n3176), .B1(n2732), .B2(n2944), .ZN(n2595)
         );
  AOI221_X1 U2942 ( .B1(n2949), .B2(n2900), .C1(n2947), .C2(n3323), .A(n2597), 
        .ZN(n2596) );
  OAI211_X1 U2943 ( .C1(n2942), .C2(n822), .A(n2592), .B(n2593), .ZN(n1017) );
  AOI22_X1 U2944 ( .A1(n2946), .A2(n3174), .B1(n2731), .B2(n2944), .ZN(n2592)
         );
  AOI221_X1 U2945 ( .B1(n2949), .B2(n2902), .C1(n2947), .C2(n3324), .A(n2594), 
        .ZN(n2593) );
  OAI211_X1 U2946 ( .C1(n2941), .C2(n817), .A(n2577), .B(n2578), .ZN(n1022) );
  AOI22_X1 U2947 ( .A1(n2946), .A2(n3164), .B1(n2726), .B2(n2944), .ZN(n2577)
         );
  AOI221_X1 U2948 ( .B1(n2508), .B2(n2895), .C1(n2947), .C2(n3329), .A(n2579), 
        .ZN(n2578) );
  OAI211_X1 U2949 ( .C1(n3112), .C2(n816), .A(n2574), .B(n2575), .ZN(n1023) );
  AOI22_X1 U2950 ( .A1(n2946), .A2(n3162), .B1(n2725), .B2(n2944), .ZN(n2574)
         );
  AOI221_X1 U2951 ( .B1(n2508), .B2(n2905), .C1(n2947), .C2(n3330), .A(n2576), 
        .ZN(n2575) );
  OAI211_X1 U2952 ( .C1(n2941), .C2(n815), .A(n2571), .B(n2572), .ZN(n1024) );
  AOI22_X1 U2953 ( .A1(n2946), .A2(n3160), .B1(n2724), .B2(n2944), .ZN(n2571)
         );
  AOI221_X1 U2954 ( .B1(n2508), .B2(n2897), .C1(n2947), .C2(n3331), .A(n2573), 
        .ZN(n2572) );
  OAI211_X1 U2955 ( .C1(n3112), .C2(n814), .A(n2568), .B(n2569), .ZN(n1025) );
  AOI22_X1 U2956 ( .A1(n2946), .A2(n3158), .B1(n2723), .B2(n2944), .ZN(n2568)
         );
  AOI221_X1 U2957 ( .B1(n2508), .B2(n2845), .C1(n2947), .C2(n3332), .A(n2570), 
        .ZN(n2569) );
  OAI211_X1 U2958 ( .C1(n2942), .C2(n1350), .A(n2612), .B(n2613), .ZN(n1011)
         );
  AOI221_X1 U2959 ( .B1(n2511), .B2(n3318), .C1(n2949), .C2(n2893), .A(n2611), 
        .ZN(n2613) );
  AOI22_X1 U2960 ( .A1(n2946), .A2(n3193), .B1(n2944), .B2(n2770), .ZN(n2612)
         );
  OAI211_X1 U2961 ( .C1(n3112), .C2(n813), .A(n2565), .B(n2566), .ZN(n1026) );
  AOI221_X1 U2962 ( .B1(n2949), .B2(n2871), .C1(n2947), .C2(n3333), .A(n2567), 
        .ZN(n2566) );
  AOI22_X1 U2963 ( .A1(n2512), .A2(n3156), .B1(n2722), .B2(n2943), .ZN(n2565)
         );
  OAI22_X1 U2964 ( .A1(nq[16]), .A2(n2945), .B1(nqp1[16]), .B2(n2510), .ZN(
        n2567) );
  OAI211_X1 U2965 ( .C1(n2942), .C2(n812), .A(n2562), .B(n2563), .ZN(n1027) );
  AOI221_X1 U2966 ( .B1(n2949), .B2(n2877), .C1(n2947), .C2(n3334), .A(n2564), 
        .ZN(n2563) );
  AOI22_X1 U2967 ( .A1(n2512), .A2(n3154), .B1(n2721), .B2(n2943), .ZN(n2562)
         );
  OAI22_X1 U2968 ( .A1(nq[15]), .A2(n2945), .B1(nqp1[15]), .B2(n2510), .ZN(
        n2564) );
  OAI211_X1 U2969 ( .C1(n3112), .C2(n811), .A(n2559), .B(n2560), .ZN(n1028) );
  AOI221_X1 U2970 ( .B1(n2949), .B2(n2823), .C1(n2947), .C2(n3335), .A(n2561), 
        .ZN(n2560) );
  AOI22_X1 U2971 ( .A1(n2512), .A2(n3152), .B1(n2720), .B2(n2943), .ZN(n2559)
         );
  OAI22_X1 U2972 ( .A1(nq[14]), .A2(n2945), .B1(nqp1[14]), .B2(n2510), .ZN(
        n2561) );
  OAI211_X1 U2973 ( .C1(n3112), .C2(n810), .A(n2556), .B(n2557), .ZN(n1029) );
  AOI221_X1 U2974 ( .B1(n2949), .B2(n2821), .C1(n2947), .C2(n3336), .A(n2558), 
        .ZN(n2557) );
  AOI22_X1 U2975 ( .A1(n2512), .A2(n3150), .B1(n2719), .B2(n2943), .ZN(n2556)
         );
  OAI22_X1 U2976 ( .A1(nq[13]), .A2(n2945), .B1(nqp1[13]), .B2(n2510), .ZN(
        n2558) );
  OAI211_X1 U2977 ( .C1(n2941), .C2(n809), .A(n2553), .B(n2554), .ZN(n1030) );
  AOI221_X1 U2978 ( .B1(n2949), .B2(n2819), .C1(n2947), .C2(n3337), .A(n2555), 
        .ZN(n2554) );
  AOI22_X1 U2979 ( .A1(n2946), .A2(n3148), .B1(n2718), .B2(n2943), .ZN(n2553)
         );
  OAI22_X1 U2980 ( .A1(nq[12]), .A2(n2945), .B1(nqp1[12]), .B2(n2510), .ZN(
        n2555) );
  OAI211_X1 U2981 ( .C1(n3112), .C2(n808), .A(n2550), .B(n2551), .ZN(n1031) );
  AOI221_X1 U2982 ( .B1(n2949), .B2(n2873), .C1(n2947), .C2(n3338), .A(n2552), 
        .ZN(n2551) );
  AOI22_X1 U2983 ( .A1(n2512), .A2(n3146), .B1(n2717), .B2(n2943), .ZN(n2550)
         );
  OAI22_X1 U2984 ( .A1(nq[11]), .A2(n2945), .B1(nqp1[11]), .B2(n2948), .ZN(
        n2552) );
  OAI211_X1 U2985 ( .C1(n3112), .C2(n807), .A(n2547), .B(n2548), .ZN(n1032) );
  AOI221_X1 U2986 ( .B1(n2949), .B2(n2817), .C1(n2947), .C2(n3339), .A(n2549), 
        .ZN(n2548) );
  AOI22_X1 U2987 ( .A1(n2512), .A2(n3144), .B1(n2716), .B2(n2943), .ZN(n2547)
         );
  OAI22_X1 U2988 ( .A1(nq[10]), .A2(n2945), .B1(nqp1[10]), .B2(n2948), .ZN(
        n2549) );
  OAI211_X1 U2989 ( .C1(n3112), .C2(n806), .A(n2544), .B(n2545), .ZN(n1033) );
  AOI221_X1 U2990 ( .B1(n2949), .B2(n2851), .C1(n2947), .C2(n3340), .A(n2546), 
        .ZN(n2545) );
  AOI22_X1 U2991 ( .A1(n2512), .A2(n3142), .B1(n2715), .B2(n2943), .ZN(n2544)
         );
  OAI22_X1 U2992 ( .A1(nq[9]), .A2(n2945), .B1(nqp1[9]), .B2(n2948), .ZN(n2546) );
  OAI211_X1 U2993 ( .C1(n2941), .C2(n805), .A(n2541), .B(n2542), .ZN(n1034) );
  AOI221_X1 U2994 ( .B1(n2949), .B2(n2854), .C1(n2947), .C2(n3341), .A(n2543), 
        .ZN(n2542) );
  AOI22_X1 U2995 ( .A1(n2946), .A2(n3140), .B1(n2714), .B2(n2943), .ZN(n2541)
         );
  OAI22_X1 U2996 ( .A1(nq[8]), .A2(n2945), .B1(nqp1[8]), .B2(n2948), .ZN(n2543) );
  OAI211_X1 U2997 ( .C1(n3112), .C2(n804), .A(n2538), .B(n2539), .ZN(n1035) );
  AOI221_X1 U2998 ( .B1(n2949), .B2(n2859), .C1(n2511), .C2(n3342), .A(n2540), 
        .ZN(n2539) );
  AOI22_X1 U2999 ( .A1(n2946), .A2(n3138), .B1(n2713), .B2(n2943), .ZN(n2538)
         );
  OAI22_X1 U3000 ( .A1(nq[7]), .A2(n2945), .B1(nqp1[7]), .B2(n2948), .ZN(n2540) );
  OAI211_X1 U3001 ( .C1(n2941), .C2(n803), .A(n2535), .B(n2536), .ZN(n1036) );
  AOI221_X1 U3002 ( .B1(n2949), .B2(n2862), .C1(n2511), .C2(n3343), .A(n2537), 
        .ZN(n2536) );
  AOI22_X1 U3003 ( .A1(n2946), .A2(n3136), .B1(n2712), .B2(n2943), .ZN(n2535)
         );
  OAI22_X1 U3004 ( .A1(nq[6]), .A2(n2945), .B1(nqp1[6]), .B2(n2948), .ZN(n2537) );
  OAI211_X1 U3005 ( .C1(n3112), .C2(n802), .A(n2532), .B(n2533), .ZN(n1037) );
  AOI221_X1 U3006 ( .B1(n2949), .B2(n2837), .C1(n2511), .C2(n3344), .A(n2534), 
        .ZN(n2533) );
  AOI22_X1 U3007 ( .A1(n2946), .A2(n3134), .B1(n2711), .B2(n2943), .ZN(n2532)
         );
  OAI22_X1 U3008 ( .A1(nq[5]), .A2(n2945), .B1(nqp1[5]), .B2(n2948), .ZN(n2534) );
  NAND2_X1 U3009 ( .A1(n2616), .A2(n2617), .ZN(n2615) );
  NOR4_X1 U3010 ( .A1(n2622), .A2(n2623), .A3(n2624), .A4(n2625), .ZN(n2616)
         );
  NOR4_X1 U3011 ( .A1(n2618), .A2(n2619), .A3(n2620), .A4(n2621), .ZN(n2617)
         );
  NAND4_X1 U3012 ( .A1(n2749), .A2(n2750), .A3(n2751), .A4(n2752), .ZN(n2622)
         );
  AOI221_X1 U3013 ( .B1(n2925), .B2(n3285), .C1(n2508), .C2(n2891), .A(n2509), 
        .ZN(n2507) );
  AOI221_X1 U3014 ( .B1(n2511), .B2(n3349), .C1(n2946), .C2(n3187), .A(n2513), 
        .ZN(n2506) );
  OAI22_X1 U3015 ( .A1(nqp1[0]), .A2(n2948), .B1(n3192), .B2(n2347), .ZN(n2509) );
  AOI221_X1 U3016 ( .B1(n2925), .B2(n3281), .C1(n2508), .C2(n2868), .A(n2528), 
        .ZN(n2527) );
  AOI221_X1 U3017 ( .B1(n2511), .B2(n3345), .C1(n2946), .C2(n3131), .A(n2530), 
        .ZN(n2526) );
  AOI221_X1 U3018 ( .B1(n2925), .B2(n3282), .C1(n2508), .C2(n2865), .A(n2524), 
        .ZN(n2523) );
  AOI221_X1 U3019 ( .B1(n2511), .B2(n3346), .C1(n2946), .C2(n3128), .A(n2525), 
        .ZN(n2522) );
  OAI22_X1 U3020 ( .A1(nqp1[3]), .A2(n2948), .B1(n3189), .B2(n2347), .ZN(n2524) );
  AOI221_X1 U3021 ( .B1(n2925), .B2(n3283), .C1(n2508), .C2(n2878), .A(n2520), 
        .ZN(n2519) );
  AOI221_X1 U3022 ( .B1(n2511), .B2(n3347), .C1(n2946), .C2(n3125), .A(n2521), 
        .ZN(n2518) );
  OAI22_X1 U3023 ( .A1(nqp1[2]), .A2(n2948), .B1(n3190), .B2(n2347), .ZN(n2520) );
  AOI221_X1 U3024 ( .B1(n2925), .B2(n3284), .C1(n2508), .C2(n2903), .A(n2516), 
        .ZN(n2515) );
  AOI221_X1 U3025 ( .B1(n2511), .B2(n3348), .C1(n2946), .C2(n3122), .A(n2517), 
        .ZN(n2514) );
  OAI22_X1 U3026 ( .A1(nqp1[1]), .A2(n2948), .B1(n3191), .B2(n2347), .ZN(n2516) );
  AND2_X1 U3027 ( .A1(n941), .A2(n2929), .ZN(n2502) );
  INV_X1 U3028 ( .A(n2346), .ZN(n3028) );
  AOI22_X1 U3029 ( .A1(n2974), .A2(sdata_o[31]), .B1(n2971), .B2(n1829), .ZN(
        n2346) );
  OR2_X1 U3030 ( .A1(n2769), .A2(n2366), .ZN(n2347) );
  NOR3_X1 U3031 ( .A1(n3110), .A2(n934), .A3(n2408), .ZN(n2318) );
  OAI211_X1 U3032 ( .C1(n941), .C2(n2941), .A(n2940), .B(n3100), .ZN(n1293) );
  OAI22_X1 U3033 ( .A1(n2402), .A2(n2638), .B1(n2958), .B2(n3222), .ZN(n1261)
         );
  OAI22_X1 U3034 ( .A1(n2960), .A2(n2639), .B1(n2958), .B2(n3221), .ZN(n1260)
         );
  OAI22_X1 U3035 ( .A1(n2402), .A2(n2640), .B1(n2958), .B2(n3207), .ZN(n1259)
         );
  OAI22_X1 U3036 ( .A1(n2960), .A2(n2637), .B1(n2959), .B2(n3223), .ZN(n1262)
         );
  OAI22_X1 U3037 ( .A1(n2770), .A2(n2957), .B1(n3058), .B2(n2953), .ZN(n1124)
         );
  OAI22_X1 U3038 ( .A1(n2703), .A2(n2955), .B1(n3115), .B2(n2954), .ZN(n1155)
         );
  OAI22_X1 U3039 ( .A1(n2713), .A2(n2955), .B1(n3137), .B2(n2954), .ZN(n1148)
         );
  OAI22_X1 U3040 ( .A1(n2712), .A2(n2955), .B1(n3135), .B2(n2954), .ZN(n1149)
         );
  OAI22_X1 U3041 ( .A1(n2711), .A2(n2955), .B1(n3133), .B2(n2954), .ZN(n1150)
         );
  OAI22_X1 U3042 ( .A1(n2710), .A2(n2955), .B1(n3130), .B2(n2954), .ZN(n1151)
         );
  OAI22_X1 U3043 ( .A1(n2709), .A2(n2956), .B1(n3127), .B2(n2954), .ZN(n1152)
         );
  OAI22_X1 U3044 ( .A1(n2707), .A2(n2955), .B1(n3124), .B2(n2954), .ZN(n1153)
         );
  OAI22_X1 U3045 ( .A1(n2705), .A2(n2956), .B1(n3121), .B2(n2954), .ZN(n1154)
         );
  OAI22_X1 U3046 ( .A1(n2768), .A2(n2406), .B1(n2940), .B2(n3286), .ZN(n1227)
         );
  OAI22_X1 U3047 ( .A1(n2736), .A2(n2957), .B1(n3183), .B2(n2953), .ZN(n1125)
         );
  OAI22_X1 U3048 ( .A1(n2735), .A2(n2957), .B1(n3181), .B2(n2953), .ZN(n1126)
         );
  OAI22_X1 U3049 ( .A1(n2734), .A2(n2957), .B1(n3179), .B2(n2953), .ZN(n1127)
         );
  OAI22_X1 U3050 ( .A1(n2733), .A2(n2955), .B1(n3177), .B2(n2953), .ZN(n1128)
         );
  OAI22_X1 U3051 ( .A1(n2732), .A2(n2955), .B1(n3175), .B2(n2953), .ZN(n1129)
         );
  OAI22_X1 U3052 ( .A1(n2731), .A2(n2956), .B1(n3173), .B2(n2953), .ZN(n1130)
         );
  OAI22_X1 U3053 ( .A1(n2730), .A2(n2955), .B1(n3171), .B2(n2953), .ZN(n1131)
         );
  OAI22_X1 U3054 ( .A1(n2729), .A2(n2955), .B1(n3169), .B2(n2953), .ZN(n1132)
         );
  OAI22_X1 U3055 ( .A1(n2728), .A2(n2956), .B1(n3167), .B2(n2953), .ZN(n1133)
         );
  OAI22_X1 U3056 ( .A1(n2727), .A2(n2955), .B1(n3165), .B2(n2953), .ZN(n1134)
         );
  OAI22_X1 U3057 ( .A1(n2726), .A2(n2956), .B1(n3163), .B2(n2953), .ZN(n1135)
         );
  OAI22_X1 U3058 ( .A1(n2725), .A2(n2955), .B1(n3161), .B2(n2954), .ZN(n1136)
         );
  OAI22_X1 U3059 ( .A1(n2724), .A2(n2956), .B1(n3159), .B2(n2954), .ZN(n1137)
         );
  OAI22_X1 U3060 ( .A1(n2723), .A2(n2955), .B1(n3157), .B2(n2954), .ZN(n1138)
         );
  OAI22_X1 U3061 ( .A1(n2722), .A2(n2956), .B1(n3155), .B2(n2954), .ZN(n1139)
         );
  OAI22_X1 U3062 ( .A1(n2721), .A2(n2955), .B1(n3153), .B2(n2954), .ZN(n1140)
         );
  OAI22_X1 U3063 ( .A1(n2720), .A2(n2955), .B1(n3151), .B2(n2954), .ZN(n1141)
         );
  OAI22_X1 U3064 ( .A1(n2719), .A2(n2955), .B1(n3149), .B2(n2954), .ZN(n1142)
         );
  OAI22_X1 U3065 ( .A1(n2718), .A2(n2955), .B1(n3147), .B2(n2954), .ZN(n1143)
         );
  OAI22_X1 U3066 ( .A1(n2717), .A2(n2956), .B1(n3145), .B2(n2954), .ZN(n1144)
         );
  OAI22_X1 U3067 ( .A1(n2716), .A2(n2956), .B1(n3143), .B2(n2954), .ZN(n1145)
         );
  OAI22_X1 U3068 ( .A1(n2715), .A2(n2956), .B1(n3141), .B2(n2954), .ZN(n1146)
         );
  OAI22_X1 U3069 ( .A1(n2714), .A2(n2956), .B1(n3139), .B2(n2954), .ZN(n1147)
         );
  OAI22_X1 U3070 ( .A1(n2979), .A2(n2669), .B1(n2980), .B2(n3223), .ZN(n1224)
         );
  OAI22_X1 U3071 ( .A1(n2978), .A2(n2670), .B1(n2980), .B2(n3222), .ZN(n1223)
         );
  OAI22_X1 U3072 ( .A1(n2978), .A2(n2671), .B1(n2980), .B2(n3221), .ZN(n1222)
         );
  OAI22_X1 U3073 ( .A1(n2979), .A2(n2672), .B1(n2980), .B2(n3207), .ZN(n1221)
         );
  XNOR2_X1 U3074 ( .A(n2768), .B(n1829), .ZN(n2614) );
  NAND4_X1 U3075 ( .A1(n2753), .A2(n2754), .A3(n2755), .A4(n2756), .ZN(n2621)
         );
  NAND4_X1 U3076 ( .A1(n2737), .A2(n2738), .A3(n2739), .A4(n2740), .ZN(n2625)
         );
  NAND4_X1 U3077 ( .A1(n2757), .A2(n2758), .A3(n2759), .A4(n2760), .ZN(n2620)
         );
  NAND4_X1 U3078 ( .A1(n2741), .A2(n2742), .A3(n2743), .A4(n2744), .ZN(n2624)
         );
  NAND4_X1 U3079 ( .A1(n2745), .A2(n2746), .A3(n2747), .A4(n2748), .ZN(n2623)
         );
  NAND4_X1 U3080 ( .A1(n2761), .A2(n2762), .A3(n2763), .A4(n2764), .ZN(n2619)
         );
  NAND2_X1 U3081 ( .A1(ready), .A2(i_start), .ZN(n2308) );
  INV_X1 U3082 ( .A(n2913), .ZN(n3321) );
  INV_X1 U3083 ( .A(n2813), .ZN(n3322) );
  INV_X1 U3084 ( .A(n2900), .ZN(n3323) );
  INV_X1 U3085 ( .A(n2902), .ZN(n3324) );
  INV_X1 U3086 ( .A(n2909), .ZN(n3325) );
  INV_X1 U3087 ( .A(n2911), .ZN(n3326) );
  INV_X1 U3088 ( .A(n2907), .ZN(n3327) );
  INV_X1 U3089 ( .A(n2890), .ZN(n3328) );
  INV_X1 U3090 ( .A(n2895), .ZN(n3329) );
  INV_X1 U3091 ( .A(n2905), .ZN(n3330) );
  INV_X1 U3092 ( .A(n2897), .ZN(n3331) );
  INV_X1 U3093 ( .A(n2845), .ZN(n3332) );
  INV_X1 U3094 ( .A(n2871), .ZN(n3333) );
  INV_X1 U3095 ( .A(n2877), .ZN(n3334) );
  INV_X1 U3096 ( .A(n2823), .ZN(n3335) );
  INV_X1 U3097 ( .A(n2821), .ZN(n3336) );
  INV_X1 U3098 ( .A(n2819), .ZN(n3337) );
  INV_X1 U3099 ( .A(n2873), .ZN(n3338) );
  INV_X1 U3100 ( .A(n2851), .ZN(n3340) );
  INV_X1 U3101 ( .A(n2854), .ZN(n3341) );
  INV_X1 U3102 ( .A(n2859), .ZN(n3342) );
  INV_X1 U3103 ( .A(n2862), .ZN(n3343) );
  INV_X1 U3104 ( .A(n2837), .ZN(n3344) );
  INV_X1 U3105 ( .A(n2916), .ZN(n3286) );
  INV_X1 U3106 ( .A(n2893), .ZN(n3318) );
  INV_X1 U3107 ( .A(n2891), .ZN(n3349) );
  INV_X1 U3108 ( .A(n2868), .ZN(n3345) );
  INV_X1 U3109 ( .A(n2865), .ZN(n3346) );
  INV_X1 U3110 ( .A(n2878), .ZN(n3347) );
  OAI22_X1 U3111 ( .A1(n2453), .A2(n3110), .B1(n2769), .B2(n3101), .ZN(n1113)
         );
  INV_X1 U3112 ( .A(n2453), .ZN(n3101) );
  NOR2_X1 U3113 ( .A1(n2973), .A2(n2320), .ZN(n2453) );
  INV_X1 U3114 ( .A(n2817), .ZN(n3339) );
  INV_X1 U3115 ( .A(n2903), .ZN(n3348) );
  BUF_X1 U3116 ( .A(i_rst), .Z(n3019) );
  BUF_X1 U3117 ( .A(i_rst), .Z(n3020) );
  OAI211_X1 U3118 ( .C1(n2942), .C2(n825), .A(n2601), .B(n2602), .ZN(n1014) );
  OAI22_X1 U3119 ( .A1(n2458), .A2(n3284), .B1(n3088), .B2(n2457), .ZN(n1104)
         );
  AND2_X1 U3120 ( .A1(n2949), .A2(i_divisor[29]), .ZN(n2932) );
  AND2_X1 U3121 ( .A1(n2511), .A2(n3320), .ZN(n2933) );
  NOR3_X1 U3122 ( .A1(n2932), .A2(n2933), .A3(n2606), .ZN(n2605) );
  INV_X1 U3123 ( .A(n2841), .ZN(n3320) );
  OR2_X1 U3124 ( .A1(n2761), .A2(n2975), .ZN(n2934) );
  OR2_X1 U3125 ( .A1(n2941), .A2(n701), .ZN(n2935) );
  AND2_X1 U3126 ( .A1(n2968), .A2(PR_1[30]), .ZN(n2936) );
  AND2_X1 U3127 ( .A1(q[30]), .A2(n2356), .ZN(n2937) );
  INV_X1 U3128 ( .A(n2976), .ZN(n2975) );
  INV_X1 U3129 ( .A(n2928), .ZN(n2968) );
  AOI22_X1 U3130 ( .A1(q[1]), .A2(n2356), .B1(qp1[1]), .B2(n2357), .ZN(n2367)
         );
  OAI221_X1 U3131 ( .B1(n2358), .B2(n3348), .C1(n2964), .C2(n3121), .A(n2421), 
        .ZN(n1185) );
  NAND2_X1 U3132 ( .A1(shifted_o[3]), .A2(n3103), .ZN(n2418) );
  NOR2_X1 U3133 ( .A1(n2609), .A2(n2789), .ZN(n2608) );
  OAI22_X1 U3134 ( .A1(n2456), .A2(n3285), .B1(n3089), .B2(n2457), .ZN(n1105)
         );
  OAI22_X1 U3135 ( .A1(nq[29]), .A2(n2945), .B1(nqp1[29]), .B2(n2510), .ZN(
        n2606) );
  OAI211_X1 U3136 ( .C1(n2942), .C2(n826), .A(n2604), .B(n2605), .ZN(n1013) );
  AOI22_X1 U3137 ( .A1(q[0]), .A2(n2356), .B1(qp1[0]), .B2(n2357), .ZN(n2364)
         );
  AND2_X1 U3138 ( .A1(n2949), .A2(i_divisor[30]), .ZN(n2938) );
  AND2_X1 U3139 ( .A1(n2511), .A2(n3319), .ZN(n2939) );
  OAI221_X1 U3140 ( .B1(n2358), .B2(n3339), .C1(n2964), .C2(n3143), .A(n2430), 
        .ZN(n1176) );
  INV_X1 U3141 ( .A(n2927), .ZN(n2943) );
  INV_X1 U3142 ( .A(n2927), .ZN(n2944) );
  INV_X1 U3143 ( .A(n2925), .ZN(n2945) );
  INV_X1 U3144 ( .A(n2344), .ZN(n2976) );
  CLKBUF_X1 U3145 ( .A(n3018), .Z(n2984) );
  CLKBUF_X1 U3146 ( .A(n3018), .Z(n2985) );
  CLKBUF_X1 U3147 ( .A(n3018), .Z(n2986) );
  CLKBUF_X1 U3148 ( .A(n3018), .Z(n2987) );
  CLKBUF_X1 U3149 ( .A(n3018), .Z(n2988) );
  CLKBUF_X1 U3150 ( .A(n3018), .Z(n2989) );
  CLKBUF_X1 U3151 ( .A(n3017), .Z(n2990) );
  CLKBUF_X1 U3152 ( .A(n3017), .Z(n2991) );
  CLKBUF_X1 U3153 ( .A(n3017), .Z(n2992) );
  CLKBUF_X1 U3154 ( .A(n3017), .Z(n2993) );
  CLKBUF_X1 U3155 ( .A(n3017), .Z(n2994) );
  CLKBUF_X1 U3156 ( .A(n3017), .Z(n2995) );
  CLKBUF_X1 U3157 ( .A(n3016), .Z(n2996) );
  CLKBUF_X1 U3158 ( .A(n3016), .Z(n2997) );
  CLKBUF_X1 U3159 ( .A(n3016), .Z(n2998) );
  CLKBUF_X1 U3160 ( .A(n3016), .Z(n2999) );
  CLKBUF_X1 U3161 ( .A(n3016), .Z(n3000) );
  CLKBUF_X1 U3162 ( .A(n3016), .Z(n3001) );
  CLKBUF_X1 U3163 ( .A(n3015), .Z(n3002) );
  CLKBUF_X1 U3164 ( .A(n3015), .Z(n3003) );
  CLKBUF_X1 U3165 ( .A(n3015), .Z(n3004) );
  CLKBUF_X1 U3166 ( .A(n3015), .Z(n3005) );
  CLKBUF_X1 U3167 ( .A(n3015), .Z(n3006) );
  CLKBUF_X1 U3168 ( .A(n3015), .Z(n3007) );
  CLKBUF_X1 U3169 ( .A(n3014), .Z(n3008) );
  CLKBUF_X1 U3170 ( .A(n3014), .Z(n3009) );
  CLKBUF_X1 U3171 ( .A(n3014), .Z(n3010) );
  CLKBUF_X1 U3172 ( .A(n3014), .Z(n3011) );
  CLKBUF_X1 U3173 ( .A(n3014), .Z(n3012) );
  CLKBUF_X1 U3174 ( .A(n3014), .Z(n3013) );
  OAI22_X1 \shifter_0/U31  ( .A1(\shifter_0/n13 ), .A2(\shifter_0/n6 ), .B1(
        \shifter_0/n21 ), .B2(\shifter_0/n7 ), .ZN(\shifter_0/n9 ) );
  OAI22_X1 \shifter_0/U30  ( .A1(\shifter_0/n32 ), .A2(\shifter_0/n8 ), .B1(
        shifted_o[3]), .B2(\shifter_0/n7 ), .ZN(shifted_o[1]) );
  OAI22_X1 \shifter_0/U28  ( .A1(\shifter_0/n31 ), .A2(\shifter_0/n6 ), .B1(
        shifted_o[3]), .B2(\shifter_0/n7 ), .ZN(shifted_o[2]) );
  OAI22_X1 \shifter_0/U27  ( .A1(\shifter_0/n9 ), .A2(\shifter_0/n10 ), .B1(
        shifted_o[3]), .B2(\shifter_0/n11 ), .ZN(shifted_o[0]) );
  XNOR2_X1 \shifter_0/U26  ( .A(sdata[31]), .B(sdata[22]), .ZN(\shifter_0/n14 ) );
  XNOR2_X1 \shifter_0/U25  ( .A(sdata[31]), .B(sdata[24]), .ZN(\shifter_0/n16 ) );
  NAND2_X1 \shifter_0/U24  ( .A1(\shifter_0/n16 ), .A2(\shifter_0/n31 ), .ZN(
        \shifter_0/n11 ) );
  XNOR2_X1 \shifter_0/U23  ( .A(sdata[31]), .B(sdata[27]), .ZN(\shifter_0/n18 ) );
  XOR2_X1 \shifter_0/U22  ( .A(sdata[31]), .B(sdata[23]), .Z(\shifter_0/n30 )
         );
  NOR2_X1 \shifter_0/U21  ( .A1(\shifter_0/n30 ), .A2(\shifter_0/n11 ), .ZN(
        shifted_o[3]) );
  XNOR2_X1 \shifter_0/U20  ( .A(sdata[31]), .B(sdata[25]), .ZN(\shifter_0/n17 ) );
  INV_X1 \shifter_0/U19  ( .A(\shifter_0/n8 ), .ZN(\shifter_0/n4 ) );
  XNOR2_X1 \shifter_0/U18  ( .A(sdata[31]), .B(sdata[26]), .ZN(\shifter_0/n13 ) );
  XNOR2_X1 \shifter_0/U17  ( .A(sdata[31]), .B(sdata[28]), .ZN(\shifter_0/n19 ) );
  INV_X1 \shifter_0/U16  ( .A(\shifter_0/n11 ), .ZN(\shifter_0/n1 ) );
  XNOR2_X1 \shifter_0/U15  ( .A(sdata[31]), .B(sdata[30]), .ZN(\shifter_0/n20 ) );
  INV_X1 \shifter_0/U14  ( .A(\shifter_0/n6 ), .ZN(\shifter_0/n32 ) );
  INV_X1 \shifter_0/U13  ( .A(\shifter_0/n7 ), .ZN(\shifter_0/n31 ) );
  OAI21_X1 \shifter_0/U12  ( .B1(\shifter_0/n25 ), .B2(\shifter_0/n12 ), .A(
        \shifter_0/n20 ), .ZN(\shifter_0/n10 ) );
  INV_X1 \shifter_0/U11  ( .A(\shifter_0/n12 ), .ZN(\shifter_0/n33 ) );
  NAND2_X1 \shifter_0/U10  ( .A1(\shifter_0/n33 ), .A2(\shifter_0/n20 ), .ZN(
        \shifter_0/n8 ) );
  AND3_X1 \shifter_0/U9  ( .A1(\shifter_0/n19 ), .A2(\shifter_0/n20 ), .A3(
        \shifter_0/n33 ), .ZN(\shifter_0/n25 ) );
  AND2_X1 \shifter_0/U8  ( .A1(\shifter_0/n32 ), .A2(\shifter_0/n13 ), .ZN(
        \shifter_0/n24 ) );
  NAND2_X1 \shifter_0/U7  ( .A1(\shifter_0/n18 ), .A2(\shifter_0/n25 ), .ZN(
        \shifter_0/n6 ) );
  NAND2_X1 \shifter_0/U6  ( .A1(\shifter_0/n17 ), .A2(\shifter_0/n24 ), .ZN(
        \shifter_0/n7 ) );
  AND2_X1 \shifter_0/U5  ( .A1(\shifter_0/n14 ), .A2(shifted_o[3]), .ZN(
        \shifter_0/n21 ) );
  INV_X1 \shifter_0/U3  ( .A(1'b1), .ZN(\shifter_0/o_shifted[4] ) );
  XOR2_X1 \shifter_0/U29  ( .A(sdata[31]), .B(sdata[29]), .Z(\shifter_0/n12 )
         );
  AOI22_X1 \shifter_0/shift_1b_0/U70  ( .A1(\shifter_0/shift_1b_0/n65 ), .A2(
        sdata[9]), .B1(sdata[8]), .B2(\shifter_0/shift_1b_0/n69 ), .ZN(
        \shifter_0/shift_1b_0/n33 ) );
  INV_X1 \shifter_0/shift_1b_0/U69  ( .A(\shifter_0/shift_1b_0/n33 ), .ZN(
        \shifter_0/data_1 [9]) );
  AND2_X1 \shifter_0/shift_1b_0/U68  ( .A1(\shifter_0/shift_1b_0/n65 ), .A2(
        sdata[0]), .ZN(\shifter_0/data_1 [0]) );
  AOI22_X1 \shifter_0/shift_1b_0/U67  ( .A1(\shifter_0/shift_1b_0/n68 ), .A2(
        sdata[9]), .B1(\shifter_0/shift_1b_0/n66 ), .B2(sdata[10]), .ZN(
        \shifter_0/shift_1b_0/n63 ) );
  INV_X1 \shifter_0/shift_1b_0/U66  ( .A(\shifter_0/shift_1b_0/n63 ), .ZN(
        \shifter_0/data_1 [10]) );
  AOI22_X1 \shifter_0/shift_1b_0/U65  ( .A1(\shifter_0/shift_1b_0/n65 ), .A2(
        sdata[11]), .B1(\shifter_0/shift_1b_0/n69 ), .B2(sdata[10]), .ZN(
        \shifter_0/shift_1b_0/n62 ) );
  INV_X1 \shifter_0/shift_1b_0/U64  ( .A(\shifter_0/shift_1b_0/n62 ), .ZN(
        \shifter_0/data_1 [11]) );
  AOI22_X1 \shifter_0/shift_1b_0/U63  ( .A1(\shifter_0/shift_1b_0/n66 ), .A2(
        sdata[1]), .B1(\shifter_0/shift_1b_0/n68 ), .B2(sdata[0]), .ZN(
        \shifter_0/shift_1b_0/n53 ) );
  INV_X1 \shifter_0/shift_1b_0/U62  ( .A(\shifter_0/shift_1b_0/n53 ), .ZN(
        \shifter_0/data_1 [1]) );
  AOI22_X1 \shifter_0/shift_1b_0/U61  ( .A1(\shifter_0/shift_1b_0/n65 ), .A2(
        sdata[2]), .B1(\shifter_0/shift_1b_0/n67 ), .B2(sdata[1]), .ZN(
        \shifter_0/shift_1b_0/n42 ) );
  INV_X1 \shifter_0/shift_1b_0/U60  ( .A(\shifter_0/shift_1b_0/n42 ), .ZN(
        \shifter_0/data_1 [2]) );
  AOI22_X1 \shifter_0/shift_1b_0/U59  ( .A1(\shifter_0/shift_1b_0/n66 ), .A2(
        sdata[21]), .B1(\shifter_0/n20 ), .B2(sdata[20]), .ZN(
        \shifter_0/shift_1b_0/n51 ) );
  INV_X1 \shifter_0/shift_1b_0/U58  ( .A(\shifter_0/shift_1b_0/n51 ), .ZN(
        \shifter_0/data_1 [21]) );
  AOI22_X1 \shifter_0/shift_1b_0/U57  ( .A1(\shifter_0/shift_1b_0/n66 ), .A2(
        sdata[20]), .B1(\shifter_0/n20 ), .B2(sdata[19]), .ZN(
        \shifter_0/shift_1b_0/n52 ) );
  INV_X1 \shifter_0/shift_1b_0/U56  ( .A(\shifter_0/shift_1b_0/n52 ), .ZN(
        \shifter_0/data_1 [20]) );
  AOI22_X1 \shifter_0/shift_1b_0/U55  ( .A1(\shifter_0/shift_1b_0/n66 ), .A2(
        sdata[19]), .B1(\shifter_0/n20 ), .B2(sdata[18]), .ZN(
        \shifter_0/shift_1b_0/n54 ) );
  INV_X1 \shifter_0/shift_1b_0/U54  ( .A(\shifter_0/shift_1b_0/n54 ), .ZN(
        \shifter_0/data_1 [19]) );
  AOI22_X1 \shifter_0/shift_1b_0/U53  ( .A1(\shifter_0/shift_1b_0/n66 ), .A2(
        sdata[18]), .B1(\shifter_0/n20 ), .B2(sdata[17]), .ZN(
        \shifter_0/shift_1b_0/n55 ) );
  INV_X1 \shifter_0/shift_1b_0/U52  ( .A(\shifter_0/shift_1b_0/n55 ), .ZN(
        \shifter_0/data_1 [18]) );
  AOI22_X1 \shifter_0/shift_1b_0/U51  ( .A1(\shifter_0/shift_1b_0/n65 ), .A2(
        sdata[3]), .B1(\shifter_0/shift_1b_0/n67 ), .B2(sdata[2]), .ZN(
        \shifter_0/shift_1b_0/n39 ) );
  INV_X1 \shifter_0/shift_1b_0/U50  ( .A(\shifter_0/shift_1b_0/n39 ), .ZN(
        \shifter_0/data_1 [3]) );
  AOI22_X1 \shifter_0/shift_1b_0/U49  ( .A1(\shifter_0/shift_1b_0/n65 ), .A2(
        sdata[4]), .B1(\shifter_0/shift_1b_0/n67 ), .B2(sdata[3]), .ZN(
        \shifter_0/shift_1b_0/n38 ) );
  INV_X1 \shifter_0/shift_1b_0/U48  ( .A(\shifter_0/shift_1b_0/n38 ), .ZN(
        \shifter_0/data_1 [4]) );
  AOI22_X1 \shifter_0/shift_1b_0/U47  ( .A1(\shifter_0/shift_1b_0/n65 ), .A2(
        sdata[5]), .B1(\shifter_0/shift_1b_0/n68 ), .B2(sdata[4]), .ZN(
        \shifter_0/shift_1b_0/n37 ) );
  INV_X1 \shifter_0/shift_1b_0/U46  ( .A(\shifter_0/shift_1b_0/n37 ), .ZN(
        \shifter_0/data_1 [5]) );
  AOI22_X1 \shifter_0/shift_1b_0/U45  ( .A1(\shifter_0/shift_1b_0/n65 ), .A2(
        sdata[6]), .B1(\shifter_0/shift_1b_0/n69 ), .B2(sdata[5]), .ZN(
        \shifter_0/shift_1b_0/n36 ) );
  INV_X1 \shifter_0/shift_1b_0/U44  ( .A(\shifter_0/shift_1b_0/n36 ), .ZN(
        \shifter_0/data_1 [6]) );
  AOI22_X1 \shifter_0/shift_1b_0/U43  ( .A1(\shifter_0/shift_1b_0/n65 ), .A2(
        sdata[7]), .B1(\shifter_0/shift_1b_0/n68 ), .B2(sdata[6]), .ZN(
        \shifter_0/shift_1b_0/n35 ) );
  INV_X1 \shifter_0/shift_1b_0/U42  ( .A(\shifter_0/shift_1b_0/n35 ), .ZN(
        \shifter_0/data_1 [7]) );
  AOI22_X1 \shifter_0/shift_1b_0/U41  ( .A1(\shifter_0/shift_1b_0/n65 ), .A2(
        sdata[12]), .B1(\shifter_0/shift_1b_0/n69 ), .B2(sdata[11]), .ZN(
        \shifter_0/shift_1b_0/n61 ) );
  INV_X1 \shifter_0/shift_1b_0/U40  ( .A(\shifter_0/shift_1b_0/n61 ), .ZN(
        \shifter_0/data_1 [12]) );
  AOI22_X1 \shifter_0/shift_1b_0/U39  ( .A1(\shifter_0/shift_1b_0/n65 ), .A2(
        sdata[13]), .B1(\shifter_0/shift_1b_0/n69 ), .B2(sdata[12]), .ZN(
        \shifter_0/shift_1b_0/n60 ) );
  INV_X1 \shifter_0/shift_1b_0/U38  ( .A(\shifter_0/shift_1b_0/n60 ), .ZN(
        \shifter_0/data_1 [13]) );
  AOI22_X1 \shifter_0/shift_1b_0/U37  ( .A1(\shifter_0/shift_1b_0/n66 ), .A2(
        sdata[14]), .B1(\shifter_0/shift_1b_0/n68 ), .B2(sdata[13]), .ZN(
        \shifter_0/shift_1b_0/n59 ) );
  INV_X1 \shifter_0/shift_1b_0/U36  ( .A(\shifter_0/shift_1b_0/n59 ), .ZN(
        \shifter_0/data_1 [14]) );
  AOI22_X1 \shifter_0/shift_1b_0/U35  ( .A1(\shifter_0/shift_1b_0/n65 ), .A2(
        sdata[15]), .B1(\shifter_0/shift_1b_0/n68 ), .B2(sdata[14]), .ZN(
        \shifter_0/shift_1b_0/n58 ) );
  INV_X1 \shifter_0/shift_1b_0/U34  ( .A(\shifter_0/shift_1b_0/n58 ), .ZN(
        \shifter_0/data_1 [15]) );
  AOI22_X1 \shifter_0/shift_1b_0/U33  ( .A1(\shifter_0/shift_1b_0/n66 ), .A2(
        sdata[16]), .B1(\shifter_0/shift_1b_0/n68 ), .B2(sdata[15]), .ZN(
        \shifter_0/shift_1b_0/n57 ) );
  INV_X1 \shifter_0/shift_1b_0/U32  ( .A(\shifter_0/shift_1b_0/n57 ), .ZN(
        \shifter_0/data_1 [16]) );
  AOI22_X1 \shifter_0/shift_1b_0/U31  ( .A1(\shifter_0/shift_1b_0/n66 ), .A2(
        sdata[17]), .B1(\shifter_0/shift_1b_0/n68 ), .B2(sdata[16]), .ZN(
        \shifter_0/shift_1b_0/n56 ) );
  INV_X1 \shifter_0/shift_1b_0/U30  ( .A(\shifter_0/shift_1b_0/n56 ), .ZN(
        \shifter_0/data_1 [17]) );
  AOI22_X1 \shifter_0/shift_1b_0/U29  ( .A1(\shifter_0/shift_1b_0/n66 ), .A2(
        sdata[23]), .B1(\shifter_0/shift_1b_0/n68 ), .B2(sdata[22]), .ZN(
        \shifter_0/shift_1b_0/n49 ) );
  INV_X1 \shifter_0/shift_1b_0/U28  ( .A(\shifter_0/shift_1b_0/n49 ), .ZN(
        \shifter_0/data_1 [23]) );
  AOI22_X1 \shifter_0/shift_1b_0/U27  ( .A1(\shifter_0/shift_1b_0/n66 ), .A2(
        sdata[24]), .B1(\shifter_0/n20 ), .B2(sdata[23]), .ZN(
        \shifter_0/shift_1b_0/n48 ) );
  INV_X1 \shifter_0/shift_1b_0/U26  ( .A(\shifter_0/shift_1b_0/n48 ), .ZN(
        \shifter_0/data_1 [24]) );
  AOI22_X1 \shifter_0/shift_1b_0/U25  ( .A1(\shifter_0/shift_1b_0/n66 ), .A2(
        sdata[22]), .B1(\shifter_0/shift_1b_0/n68 ), .B2(sdata[21]), .ZN(
        \shifter_0/shift_1b_0/n50 ) );
  INV_X1 \shifter_0/shift_1b_0/U24  ( .A(\shifter_0/shift_1b_0/n50 ), .ZN(
        \shifter_0/data_1 [22]) );
  AOI22_X1 \shifter_0/shift_1b_0/U23  ( .A1(\shifter_0/shift_1b_0/n65 ), .A2(
        sdata[8]), .B1(\shifter_0/shift_1b_0/n68 ), .B2(sdata[7]), .ZN(
        \shifter_0/shift_1b_0/n34 ) );
  INV_X1 \shifter_0/shift_1b_0/U22  ( .A(\shifter_0/shift_1b_0/n34 ), .ZN(
        \shifter_0/data_1 [8]) );
  AOI22_X1 \shifter_0/shift_1b_0/U21  ( .A1(\shifter_0/shift_1b_0/n65 ), .A2(
        sdata[30]), .B1(\shifter_0/shift_1b_0/n68 ), .B2(sdata[29]), .ZN(
        \shifter_0/shift_1b_0/n41 ) );
  INV_X1 \shifter_0/shift_1b_0/U20  ( .A(\shifter_0/shift_1b_0/n41 ), .ZN(
        \shifter_0/data_1 [30]) );
  AOI22_X1 \shifter_0/shift_1b_0/U19  ( .A1(\shifter_0/shift_1b_0/n66 ), .A2(
        sdata[25]), .B1(\shifter_0/shift_1b_0/n68 ), .B2(sdata[24]), .ZN(
        \shifter_0/shift_1b_0/n47 ) );
  INV_X1 \shifter_0/shift_1b_0/U18  ( .A(\shifter_0/shift_1b_0/n47 ), .ZN(
        \shifter_0/data_1 [25]) );
  AOI22_X1 \shifter_0/shift_1b_0/U17  ( .A1(\shifter_0/shift_1b_0/n66 ), .A2(
        sdata[26]), .B1(\shifter_0/shift_1b_0/n68 ), .B2(sdata[25]), .ZN(
        \shifter_0/shift_1b_0/n46 ) );
  INV_X1 \shifter_0/shift_1b_0/U16  ( .A(\shifter_0/shift_1b_0/n46 ), .ZN(
        \shifter_0/data_1 [26]) );
  AOI22_X1 \shifter_0/shift_1b_0/U15  ( .A1(\shifter_0/shift_1b_0/n66 ), .A2(
        sdata[27]), .B1(\shifter_0/shift_1b_0/n68 ), .B2(sdata[26]), .ZN(
        \shifter_0/shift_1b_0/n45 ) );
  INV_X1 \shifter_0/shift_1b_0/U14  ( .A(\shifter_0/shift_1b_0/n45 ), .ZN(
        \shifter_0/data_1 [27]) );
  AOI22_X1 \shifter_0/shift_1b_0/U13  ( .A1(\shifter_0/shift_1b_0/n65 ), .A2(
        sdata[28]), .B1(\shifter_0/shift_1b_0/n67 ), .B2(sdata[27]), .ZN(
        \shifter_0/shift_1b_0/n44 ) );
  INV_X1 \shifter_0/shift_1b_0/U12  ( .A(\shifter_0/shift_1b_0/n44 ), .ZN(
        \shifter_0/data_1 [28]) );
  AOI22_X1 \shifter_0/shift_1b_0/U11  ( .A1(\shifter_0/shift_1b_0/n65 ), .A2(
        sdata[29]), .B1(\shifter_0/shift_1b_0/n67 ), .B2(sdata[28]), .ZN(
        \shifter_0/shift_1b_0/n43 ) );
  INV_X1 \shifter_0/shift_1b_0/U10  ( .A(\shifter_0/shift_1b_0/n43 ), .ZN(
        \shifter_0/data_1 [29]) );
  AOI22_X1 \shifter_0/shift_1b_0/U9  ( .A1(\shifter_0/shift_1b_0/n65 ), .A2(
        sdata[31]), .B1(\shifter_0/shift_1b_0/n67 ), .B2(sdata[30]), .ZN(
        \shifter_0/shift_1b_0/n40 ) );
  INV_X1 \shifter_0/shift_1b_0/U8  ( .A(\shifter_0/shift_1b_0/n40 ), .ZN(
        \shifter_0/data_1 [31]) );
  BUF_X1 \shifter_0/shift_1b_0/U7  ( .A(\shifter_0/shift_1b_0/n64 ), .Z(
        \shifter_0/shift_1b_0/n69 ) );
  BUF_X1 \shifter_0/shift_1b_0/U6  ( .A(\shifter_0/shift_1b_0/n64 ), .Z(
        \shifter_0/shift_1b_0/n68 ) );
  BUF_X1 \shifter_0/shift_1b_0/U5  ( .A(\shifter_0/shift_1b_0/n69 ), .Z(
        \shifter_0/shift_1b_0/n67 ) );
  INV_X1 \shifter_0/shift_1b_0/U4  ( .A(\shifter_0/shift_1b_0/n64 ), .ZN(
        \shifter_0/shift_1b_0/n66 ) );
  INV_X1 \shifter_0/shift_1b_0/U3  ( .A(\shifter_0/n20 ), .ZN(
        \shifter_0/shift_1b_0/n65 ) );
  CLKBUF_X1 \shifter_0/shift_1b_0/U2  ( .A(\shifter_0/n20 ), .Z(
        \shifter_0/shift_1b_0/n64 ) );
  INV_X1 \shifter_0/shift_3b_0/U72  ( .A(\shifter_0/data_1 [9]), .ZN(
        \shifter_0/shift_3b_0/n39 ) );
  INV_X1 \shifter_0/shift_3b_0/U71  ( .A(\shifter_0/data_1 [0]), .ZN(
        \shifter_0/shift_3b_0/n71 ) );
  INV_X1 \shifter_0/shift_3b_0/U70  ( .A(\shifter_0/data_1 [10]), .ZN(
        \shifter_0/shift_3b_0/n70 ) );
  INV_X1 \shifter_0/shift_3b_0/U69  ( .A(\shifter_0/data_1 [11]), .ZN(
        \shifter_0/shift_3b_0/n69 ) );
  INV_X1 \shifter_0/shift_3b_0/U68  ( .A(\shifter_0/data_1 [1]), .ZN(
        \shifter_0/shift_3b_0/n54 ) );
  INV_X1 \shifter_0/shift_3b_0/U67  ( .A(\shifter_0/data_1 [2]), .ZN(
        \shifter_0/shift_3b_0/n46 ) );
  INV_X1 \shifter_0/shift_3b_0/U66  ( .A(\shifter_0/data_1 [21]), .ZN(
        \shifter_0/shift_3b_0/n52 ) );
  INV_X1 \shifter_0/shift_3b_0/U65  ( .A(\shifter_0/data_1 [20]), .ZN(
        \shifter_0/shift_3b_0/n53 ) );
  INV_X1 \shifter_0/shift_3b_0/U64  ( .A(\shifter_0/data_1 [19]), .ZN(
        \shifter_0/shift_3b_0/n55 ) );
  INV_X1 \shifter_0/shift_3b_0/U63  ( .A(\shifter_0/data_1 [18]), .ZN(
        \shifter_0/shift_3b_0/n56 ) );
  INV_X1 \shifter_0/shift_3b_0/U62  ( .A(\shifter_0/data_1 [3]), .ZN(
        \shifter_0/shift_3b_0/n45 ) );
  INV_X1 \shifter_0/shift_3b_0/U61  ( .A(\shifter_0/data_1 [4]), .ZN(
        \shifter_0/shift_3b_0/n44 ) );
  INV_X1 \shifter_0/shift_3b_0/U60  ( .A(\shifter_0/data_1 [5]), .ZN(
        \shifter_0/shift_3b_0/n43 ) );
  INV_X1 \shifter_0/shift_3b_0/U59  ( .A(\shifter_0/data_1 [6]), .ZN(
        \shifter_0/shift_3b_0/n42 ) );
  INV_X1 \shifter_0/shift_3b_0/U58  ( .A(\shifter_0/data_1 [7]), .ZN(
        \shifter_0/shift_3b_0/n41 ) );
  INV_X1 \shifter_0/shift_3b_0/U57  ( .A(\shifter_0/data_1 [12]), .ZN(
        \shifter_0/shift_3b_0/n68 ) );
  INV_X1 \shifter_0/shift_3b_0/U56  ( .A(\shifter_0/data_1 [13]), .ZN(
        \shifter_0/shift_3b_0/n67 ) );
  INV_X1 \shifter_0/shift_3b_0/U55  ( .A(\shifter_0/data_1 [14]), .ZN(
        \shifter_0/shift_3b_0/n66 ) );
  INV_X1 \shifter_0/shift_3b_0/U54  ( .A(\shifter_0/data_1 [15]), .ZN(
        \shifter_0/shift_3b_0/n59 ) );
  INV_X1 \shifter_0/shift_3b_0/U53  ( .A(\shifter_0/data_1 [16]), .ZN(
        \shifter_0/shift_3b_0/n58 ) );
  INV_X1 \shifter_0/shift_3b_0/U52  ( .A(\shifter_0/data_1 [17]), .ZN(
        \shifter_0/shift_3b_0/n57 ) );
  INV_X1 \shifter_0/shift_3b_0/U51  ( .A(\shifter_0/data_1 [23]), .ZN(
        \shifter_0/shift_3b_0/n50 ) );
  INV_X1 \shifter_0/shift_3b_0/U50  ( .A(\shifter_0/data_1 [24]), .ZN(
        \shifter_0/shift_3b_0/n49 ) );
  INV_X1 \shifter_0/shift_3b_0/U49  ( .A(\shifter_0/data_1 [22]), .ZN(
        \shifter_0/shift_3b_0/n51 ) );
  INV_X1 \shifter_0/shift_3b_0/U48  ( .A(\shifter_0/data_1 [8]), .ZN(
        \shifter_0/shift_3b_0/n40 ) );
  AOI22_X1 \shifter_0/shift_3b_0/U47  ( .A1(\shifter_0/shift_3b_0/n37 ), .A2(
        \shifter_0/data_1 [30]), .B1(\shifter_0/shift_3b_0/n36 ), .B2(
        \shifter_0/data_1 [28]), .ZN(\shifter_0/shift_3b_0/n65 ) );
  INV_X1 \shifter_0/shift_3b_0/U46  ( .A(\shifter_0/shift_3b_0/n65 ), .ZN(
        \shifter_0/shift_3b_0/n13 ) );
  INV_X1 \shifter_0/shift_3b_0/U45  ( .A(\shifter_0/n4 ), .ZN(
        \shifter_0/shift_3b_0/n72 ) );
  OAI21_X1 \shifter_0/shift_3b_0/U44  ( .B1(1'b0), .B2(
        \shifter_0/shift_3b_0/n72 ), .A(\shifter_0/shift_3b_0/n35 ), .ZN(
        \shifter_0/shift_3b_0/n60 ) );
  OAI21_X1 \shifter_0/shift_3b_0/U43  ( .B1(\shifter_0/shift_3b_0/n36 ), .B2(
        \shifter_0/shift_3b_0/n72 ), .A(\shifter_0/shift_3b_0/n60 ), .ZN(
        \shifter_0/shift_3b_0/shift1 ) );
  INV_X1 \shifter_0/shift_3b_0/U42  ( .A(\shifter_0/n25 ), .ZN(
        \shifter_0/shift_3b_0/n38 ) );
  AOI22_X1 \shifter_0/shift_3b_0/U41  ( .A1(\shifter_0/shift_3b_0/n37 ), .A2(
        \shifter_0/data_1 [29]), .B1(\shifter_0/shift_3b_0/n36 ), .B2(
        \shifter_0/data_1 [27]), .ZN(\shifter_0/shift_3b_0/n64 ) );
  INV_X1 \shifter_0/shift_3b_0/U40  ( .A(\shifter_0/shift_3b_0/n64 ), .ZN(
        \shifter_0/shift_3b_0/n5 ) );
  AOI22_X1 \shifter_0/shift_3b_0/U39  ( .A1(\shifter_0/shift_3b_0/n37 ), .A2(
        \shifter_0/data_1 [28]), .B1(\shifter_0/n25 ), .B2(
        \shifter_0/data_1 [26]), .ZN(\shifter_0/shift_3b_0/n63 ) );
  INV_X1 \shifter_0/shift_3b_0/U38  ( .A(\shifter_0/shift_3b_0/n63 ), .ZN(
        \shifter_0/shift_3b_0/n4 ) );
  AOI22_X1 \shifter_0/shift_3b_0/U37  ( .A1(\shifter_0/shift_3b_0/n38 ), .A2(
        \shifter_0/data_1 [27]), .B1(\shifter_0/shift_3b_0/n35 ), .B2(
        \shifter_0/data_1 [25]), .ZN(\shifter_0/shift_3b_0/n62 ) );
  INV_X1 \shifter_0/shift_3b_0/U36  ( .A(\shifter_0/shift_3b_0/n62 ), .ZN(
        \shifter_0/shift_3b_0/n3 ) );
  NOR2_X1 \shifter_0/shift_3b_0/U35  ( .A1(\shifter_0/shift_3b_0/n35 ), .A2(
        \shifter_0/shift_3b_0/n71 ), .ZN(\shifter_0/shift_3b_0/data1 [0]) );
  AOI22_X1 \shifter_0/shift_3b_0/U34  ( .A1(\shifter_0/shift_3b_0/n37 ), .A2(
        \shifter_0/data_1 [31]), .B1(\shifter_0/shift_3b_0/n36 ), .B2(
        \shifter_0/data_1 [29]), .ZN(\shifter_0/shift_3b_0/n61 ) );
  INV_X1 \shifter_0/shift_3b_0/U33  ( .A(\shifter_0/shift_3b_0/n61 ), .ZN(
        \shifter_0/shift_3b_0/n2 ) );
  NOR2_X1 \shifter_0/shift_3b_0/U32  ( .A1(\shifter_0/shift_3b_0/n35 ), .A2(
        \shifter_0/shift_3b_0/n54 ), .ZN(\shifter_0/shift_3b_0/data1 [1]) );
  OAI22_X1 \shifter_0/shift_3b_0/U31  ( .A1(\shifter_0/shift_3b_0/n36 ), .A2(
        \shifter_0/shift_3b_0/n40 ), .B1(\shifter_0/shift_3b_0/n37 ), .B2(
        \shifter_0/shift_3b_0/n42 ), .ZN(\shifter_0/shift_3b_0/n7 ) );
  OAI22_X1 \shifter_0/shift_3b_0/U30  ( .A1(\shifter_0/shift_3b_0/n35 ), .A2(
        \shifter_0/shift_3b_0/n68 ), .B1(\shifter_0/shift_3b_0/n37 ), .B2(
        \shifter_0/shift_3b_0/n70 ), .ZN(\shifter_0/shift_3b_0/n32 ) );
  OAI22_X1 \shifter_0/shift_3b_0/U29  ( .A1(\shifter_0/shift_3b_0/n36 ), .A2(
        \shifter_0/shift_3b_0/n46 ), .B1(\shifter_0/shift_3b_0/n37 ), .B2(
        \shifter_0/shift_3b_0/n71 ), .ZN(\shifter_0/shift_3b_0/n14 ) );
  INV_X1 \shifter_0/shift_3b_0/U28  ( .A(\shifter_0/data_1 [25]), .ZN(
        \shifter_0/shift_3b_0/n48 ) );
  OAI22_X1 \shifter_0/shift_3b_0/U27  ( .A1(\shifter_0/shift_3b_0/n36 ), .A2(
        \shifter_0/shift_3b_0/n48 ), .B1(\shifter_0/shift_3b_0/n37 ), .B2(
        \shifter_0/shift_3b_0/n50 ), .ZN(\shifter_0/shift_3b_0/n19 ) );
  OAI22_X1 \shifter_0/shift_3b_0/U26  ( .A1(\shifter_0/shift_3b_0/n36 ), .A2(
        \shifter_0/shift_3b_0/n50 ), .B1(\shifter_0/shift_3b_0/n38 ), .B2(
        \shifter_0/shift_3b_0/n52 ), .ZN(\shifter_0/shift_3b_0/n21 ) );
  OAI22_X1 \shifter_0/shift_3b_0/U25  ( .A1(\shifter_0/shift_3b_0/n36 ), .A2(
        \shifter_0/shift_3b_0/n51 ), .B1(\shifter_0/shift_3b_0/n38 ), .B2(
        \shifter_0/shift_3b_0/n53 ), .ZN(\shifter_0/shift_3b_0/n22 ) );
  OAI22_X1 \shifter_0/shift_3b_0/U24  ( .A1(\shifter_0/shift_3b_0/n36 ), .A2(
        \shifter_0/shift_3b_0/n52 ), .B1(\shifter_0/shift_3b_0/n38 ), .B2(
        \shifter_0/shift_3b_0/n55 ), .ZN(\shifter_0/shift_3b_0/n23 ) );
  INV_X1 \shifter_0/shift_3b_0/U23  ( .A(\shifter_0/data_1 [26]), .ZN(
        \shifter_0/shift_3b_0/n47 ) );
  OAI22_X1 \shifter_0/shift_3b_0/U22  ( .A1(\shifter_0/n25 ), .A2(
        \shifter_0/shift_3b_0/n47 ), .B1(\shifter_0/shift_3b_0/n38 ), .B2(
        \shifter_0/shift_3b_0/n49 ), .ZN(\shifter_0/shift_3b_0/n18 ) );
  OAI22_X1 \shifter_0/shift_3b_0/U21  ( .A1(\shifter_0/shift_3b_0/n36 ), .A2(
        \shifter_0/shift_3b_0/n53 ), .B1(\shifter_0/shift_3b_0/n37 ), .B2(
        \shifter_0/shift_3b_0/n56 ), .ZN(\shifter_0/shift_3b_0/n24 ) );
  OAI22_X1 \shifter_0/shift_3b_0/U20  ( .A1(\shifter_0/shift_3b_0/n36 ), .A2(
        \shifter_0/shift_3b_0/n45 ), .B1(\shifter_0/shift_3b_0/n37 ), .B2(
        \shifter_0/shift_3b_0/n54 ), .ZN(\shifter_0/shift_3b_0/n12 ) );
  OAI22_X1 \shifter_0/shift_3b_0/U19  ( .A1(\shifter_0/shift_3b_0/n36 ), .A2(
        \shifter_0/shift_3b_0/n44 ), .B1(\shifter_0/shift_3b_0/n37 ), .B2(
        \shifter_0/shift_3b_0/n46 ), .ZN(\shifter_0/shift_3b_0/n11 ) );
  OAI22_X1 \shifter_0/shift_3b_0/U18  ( .A1(\shifter_0/shift_3b_0/n35 ), .A2(
        \shifter_0/shift_3b_0/n43 ), .B1(\shifter_0/shift_3b_0/n37 ), .B2(
        \shifter_0/shift_3b_0/n45 ), .ZN(\shifter_0/shift_3b_0/n10 ) );
  OAI22_X1 \shifter_0/shift_3b_0/U17  ( .A1(\shifter_0/shift_3b_0/n35 ), .A2(
        \shifter_0/shift_3b_0/n42 ), .B1(\shifter_0/shift_3b_0/n37 ), .B2(
        \shifter_0/shift_3b_0/n44 ), .ZN(\shifter_0/shift_3b_0/n9 ) );
  OAI22_X1 \shifter_0/shift_3b_0/U16  ( .A1(\shifter_0/shift_3b_0/n35 ), .A2(
        \shifter_0/shift_3b_0/n41 ), .B1(\shifter_0/shift_3b_0/n37 ), .B2(
        \shifter_0/shift_3b_0/n43 ), .ZN(\shifter_0/shift_3b_0/n8 ) );
  OAI22_X1 \shifter_0/shift_3b_0/U15  ( .A1(\shifter_0/shift_3b_0/n35 ), .A2(
        \shifter_0/shift_3b_0/n67 ), .B1(\shifter_0/shift_3b_0/n37 ), .B2(
        \shifter_0/shift_3b_0/n69 ), .ZN(\shifter_0/shift_3b_0/n31 ) );
  OAI22_X1 \shifter_0/shift_3b_0/U14  ( .A1(\shifter_0/shift_3b_0/n35 ), .A2(
        \shifter_0/shift_3b_0/n66 ), .B1(\shifter_0/shift_3b_0/n37 ), .B2(
        \shifter_0/shift_3b_0/n68 ), .ZN(\shifter_0/shift_3b_0/n30 ) );
  OAI22_X1 \shifter_0/shift_3b_0/U13  ( .A1(\shifter_0/shift_3b_0/n36 ), .A2(
        \shifter_0/shift_3b_0/n59 ), .B1(\shifter_0/shift_3b_0/n37 ), .B2(
        \shifter_0/shift_3b_0/n67 ), .ZN(\shifter_0/shift_3b_0/n29 ) );
  OAI22_X1 \shifter_0/shift_3b_0/U12  ( .A1(\shifter_0/shift_3b_0/n36 ), .A2(
        \shifter_0/shift_3b_0/n58 ), .B1(\shifter_0/shift_3b_0/n37 ), .B2(
        \shifter_0/shift_3b_0/n66 ), .ZN(\shifter_0/shift_3b_0/n28 ) );
  OAI22_X1 \shifter_0/shift_3b_0/U11  ( .A1(\shifter_0/shift_3b_0/n36 ), .A2(
        \shifter_0/shift_3b_0/n57 ), .B1(\shifter_0/shift_3b_0/n37 ), .B2(
        \shifter_0/shift_3b_0/n59 ), .ZN(\shifter_0/shift_3b_0/n27 ) );
  OAI22_X1 \shifter_0/shift_3b_0/U10  ( .A1(\shifter_0/shift_3b_0/n36 ), .A2(
        \shifter_0/shift_3b_0/n56 ), .B1(\shifter_0/shift_3b_0/n37 ), .B2(
        \shifter_0/shift_3b_0/n58 ), .ZN(\shifter_0/shift_3b_0/n26 ) );
  OAI22_X1 \shifter_0/shift_3b_0/U9  ( .A1(\shifter_0/shift_3b_0/n36 ), .A2(
        \shifter_0/shift_3b_0/n55 ), .B1(\shifter_0/shift_3b_0/n37 ), .B2(
        \shifter_0/shift_3b_0/n57 ), .ZN(\shifter_0/shift_3b_0/n25 ) );
  OAI22_X1 \shifter_0/shift_3b_0/U8  ( .A1(\shifter_0/shift_3b_0/n36 ), .A2(
        \shifter_0/shift_3b_0/n49 ), .B1(\shifter_0/shift_3b_0/n37 ), .B2(
        \shifter_0/shift_3b_0/n51 ), .ZN(\shifter_0/shift_3b_0/n20 ) );
  OAI22_X1 \shifter_0/shift_3b_0/U7  ( .A1(\shifter_0/shift_3b_0/n37 ), .A2(
        \shifter_0/shift_3b_0/n40 ), .B1(\shifter_0/shift_3b_0/n35 ), .B2(
        \shifter_0/shift_3b_0/n70 ), .ZN(\shifter_0/shift_3b_0/n34 ) );
  OAI22_X1 \shifter_0/shift_3b_0/U6  ( .A1(\shifter_0/shift_3b_0/n35 ), .A2(
        \shifter_0/shift_3b_0/n39 ), .B1(\shifter_0/shift_3b_0/n37 ), .B2(
        \shifter_0/shift_3b_0/n41 ), .ZN(\shifter_0/shift_3b_0/n6 ) );
  OAI22_X1 \shifter_0/shift_3b_0/U5  ( .A1(\shifter_0/shift_3b_0/n37 ), .A2(
        \shifter_0/shift_3b_0/n39 ), .B1(\shifter_0/shift_3b_0/n35 ), .B2(
        \shifter_0/shift_3b_0/n69 ), .ZN(\shifter_0/shift_3b_0/n33 ) );
  BUF_X1 \shifter_0/shift_3b_0/U4  ( .A(\shifter_0/shift_3b_0/n38 ), .Z(
        \shifter_0/shift_3b_0/n37 ) );
  INV_X1 \shifter_0/shift_3b_0/U3  ( .A(\shifter_0/shift_3b_0/n38 ), .ZN(
        \shifter_0/shift_3b_0/n36 ) );
  INV_X1 \shifter_0/shift_3b_0/U2  ( .A(\shifter_0/shift_3b_0/n38 ), .ZN(
        \shifter_0/shift_3b_0/n35 ) );
  BUF_X1 \shifter_0/shift_3b_0/shift_1b_0/U68  ( .A(
        \shifter_0/shift_3b_0/shift1 ), .Z(
        \shifter_0/shift_3b_0/shift_1b_0/n64 ) );
  AOI22_X1 \shifter_0/shift_3b_0/shift_1b_0/U67  ( .A1(
        \shifter_0/shift_3b_0/shift_1b_0/n65 ), .A2(\shifter_0/shift_3b_0/n13 ), .B1(\shifter_0/shift_3b_0/shift1 ), .B2(\shifter_0/shift_3b_0/n5 ), .ZN(
        \shifter_0/shift_3b_0/shift_1b_0/n41 ) );
  INV_X1 \shifter_0/shift_3b_0/shift_1b_0/U66  ( .A(
        \shifter_0/shift_3b_0/shift_1b_0/n41 ), .ZN(\shifter_0/data_2 [30]) );
  AOI22_X1 \shifter_0/shift_3b_0/shift_1b_0/U65  ( .A1(
        \shifter_0/shift_3b_0/shift_1b_0/n65 ), .A2(\shifter_0/shift_3b_0/n2 ), 
        .B1(\shifter_0/shift_3b_0/shift_1b_0/n64 ), .B2(
        \shifter_0/shift_3b_0/n13 ), .ZN(\shifter_0/shift_3b_0/shift_1b_0/n40 ) );
  AND2_X1 \shifter_0/shift_3b_0/shift_1b_0/U64  ( .A1(
        \shifter_0/shift_3b_0/shift_1b_0/n65 ), .A2(
        \shifter_0/shift_3b_0/data1 [0]), .ZN(\shifter_0/data_2 [0]) );
  AOI22_X1 \shifter_0/shift_3b_0/shift_1b_0/U63  ( .A1(
        \shifter_0/shift_3b_0/shift_1b_0/n65 ), .A2(\shifter_0/shift_3b_0/n33 ), .B1(\shifter_0/shift_3b_0/shift_1b_0/n67 ), .B2(\shifter_0/shift_3b_0/n34 ), 
        .ZN(\shifter_0/shift_3b_0/shift_1b_0/n62 ) );
  INV_X1 \shifter_0/shift_3b_0/shift_1b_0/U62  ( .A(
        \shifter_0/shift_3b_0/shift_1b_0/n62 ), .ZN(\shifter_0/data_2 [11]) );
  AOI22_X1 \shifter_0/shift_3b_0/shift_1b_0/U61  ( .A1(
        \shifter_0/shift_3b_0/shift_1b_0/n64 ), .A2(\shifter_0/shift_3b_0/n6 ), 
        .B1(\shifter_0/shift_3b_0/shift_1b_0/n66 ), .B2(
        \shifter_0/shift_3b_0/n34 ), .ZN(\shifter_0/shift_3b_0/shift_1b_0/n63 ) );
  INV_X1 \shifter_0/shift_3b_0/shift_1b_0/U60  ( .A(
        \shifter_0/shift_3b_0/shift_1b_0/n63 ), .ZN(\shifter_0/data_2 [10]) );
  AOI22_X1 \shifter_0/shift_3b_0/shift_1b_0/U59  ( .A1(
        \shifter_0/shift_3b_0/shift_1b_0/n66 ), .A2(
        \shifter_0/shift_3b_0/data1 [1]), .B1(
        \shifter_0/shift_3b_0/shift_1b_0/n67 ), .B2(
        \shifter_0/shift_3b_0/data1 [0]), .ZN(
        \shifter_0/shift_3b_0/shift_1b_0/n53 ) );
  INV_X1 \shifter_0/shift_3b_0/shift_1b_0/U58  ( .A(
        \shifter_0/shift_3b_0/shift_1b_0/n53 ), .ZN(\shifter_0/data_2 [1]) );
  AOI22_X1 \shifter_0/shift_3b_0/shift_1b_0/U57  ( .A1(
        \shifter_0/shift_3b_0/shift_1b_0/n65 ), .A2(\shifter_0/shift_3b_0/n12 ), .B1(\shifter_0/shift_3b_0/shift_1b_0/n67 ), .B2(\shifter_0/shift_3b_0/n14 ), 
        .ZN(\shifter_0/shift_3b_0/shift_1b_0/n39 ) );
  INV_X1 \shifter_0/shift_3b_0/shift_1b_0/U56  ( .A(
        \shifter_0/shift_3b_0/shift_1b_0/n39 ), .ZN(\shifter_0/data_2 [3]) );
  AOI22_X1 \shifter_0/shift_3b_0/shift_1b_0/U55  ( .A1(
        \shifter_0/shift_3b_0/shift_1b_0/n65 ), .A2(\shifter_0/shift_3b_0/n11 ), .B1(\shifter_0/shift_3b_0/shift_1b_0/n67 ), .B2(\shifter_0/shift_3b_0/n12 ), 
        .ZN(\shifter_0/shift_3b_0/shift_1b_0/n38 ) );
  INV_X1 \shifter_0/shift_3b_0/shift_1b_0/U54  ( .A(
        \shifter_0/shift_3b_0/shift_1b_0/n38 ), .ZN(\shifter_0/data_2 [4]) );
  AOI22_X1 \shifter_0/shift_3b_0/shift_1b_0/U53  ( .A1(
        \shifter_0/shift_3b_0/shift_1b_0/n65 ), .A2(\shifter_0/shift_3b_0/n14 ), .B1(\shifter_0/shift_3b_0/shift_1b_0/n67 ), .B2(
        \shifter_0/shift_3b_0/data1 [1]), .ZN(
        \shifter_0/shift_3b_0/shift_1b_0/n42 ) );
  INV_X1 \shifter_0/shift_3b_0/shift_1b_0/U52  ( .A(
        \shifter_0/shift_3b_0/shift_1b_0/n42 ), .ZN(\shifter_0/data_2 [2]) );
  AOI22_X1 \shifter_0/shift_3b_0/shift_1b_0/U51  ( .A1(
        \shifter_0/shift_3b_0/shift_1b_0/n65 ), .A2(\shifter_0/shift_3b_0/n30 ), .B1(\shifter_0/shift_3b_0/shift_1b_0/n64 ), .B2(\shifter_0/shift_3b_0/n31 ), 
        .ZN(\shifter_0/shift_3b_0/shift_1b_0/n59 ) );
  INV_X1 \shifter_0/shift_3b_0/shift_1b_0/U50  ( .A(
        \shifter_0/shift_3b_0/shift_1b_0/n59 ), .ZN(\shifter_0/data_2 [14]) );
  AOI22_X1 \shifter_0/shift_3b_0/shift_1b_0/U49  ( .A1(
        \shifter_0/shift_3b_0/shift_1b_0/n66 ), .A2(\shifter_0/shift_3b_0/n31 ), .B1(\shifter_0/shift_3b_0/shift_1b_0/n67 ), .B2(\shifter_0/shift_3b_0/n32 ), 
        .ZN(\shifter_0/shift_3b_0/shift_1b_0/n60 ) );
  INV_X1 \shifter_0/shift_3b_0/shift_1b_0/U48  ( .A(
        \shifter_0/shift_3b_0/shift_1b_0/n60 ), .ZN(\shifter_0/data_2 [13]) );
  AOI22_X1 \shifter_0/shift_3b_0/shift_1b_0/U47  ( .A1(
        \shifter_0/shift_3b_0/shift_1b_0/n65 ), .A2(\shifter_0/shift_3b_0/n32 ), .B1(\shifter_0/shift_3b_0/shift_1b_0/n67 ), .B2(\shifter_0/shift_3b_0/n33 ), 
        .ZN(\shifter_0/shift_3b_0/shift_1b_0/n61 ) );
  INV_X1 \shifter_0/shift_3b_0/shift_1b_0/U46  ( .A(
        \shifter_0/shift_3b_0/shift_1b_0/n61 ), .ZN(\shifter_0/data_2 [12]) );
  AOI22_X1 \shifter_0/shift_3b_0/shift_1b_0/U45  ( .A1(
        \shifter_0/shift_3b_0/shift_1b_0/n65 ), .A2(\shifter_0/shift_3b_0/n8 ), 
        .B1(\shifter_0/shift_3b_0/shift_1b_0/n67 ), .B2(
        \shifter_0/shift_3b_0/n9 ), .ZN(\shifter_0/shift_3b_0/shift_1b_0/n35 )
         );
  INV_X1 \shifter_0/shift_3b_0/shift_1b_0/U44  ( .A(
        \shifter_0/shift_3b_0/shift_1b_0/n35 ), .ZN(\shifter_0/data_2 [7]) );
  AOI22_X1 \shifter_0/shift_3b_0/shift_1b_0/U43  ( .A1(
        \shifter_0/shift_3b_0/shift_1b_0/n65 ), .A2(\shifter_0/shift_3b_0/n9 ), 
        .B1(\shifter_0/shift_3b_0/shift_1b_0/n67 ), .B2(
        \shifter_0/shift_3b_0/n10 ), .ZN(\shifter_0/shift_3b_0/shift_1b_0/n36 ) );
  INV_X1 \shifter_0/shift_3b_0/shift_1b_0/U42  ( .A(
        \shifter_0/shift_3b_0/shift_1b_0/n36 ), .ZN(\shifter_0/data_2 [6]) );
  AOI22_X1 \shifter_0/shift_3b_0/shift_1b_0/U41  ( .A1(
        \shifter_0/shift_3b_0/shift_1b_0/n65 ), .A2(\shifter_0/shift_3b_0/n10 ), .B1(\shifter_0/shift_3b_0/shift_1b_0/n67 ), .B2(\shifter_0/shift_3b_0/n11 ), 
        .ZN(\shifter_0/shift_3b_0/shift_1b_0/n37 ) );
  INV_X1 \shifter_0/shift_3b_0/shift_1b_0/U40  ( .A(
        \shifter_0/shift_3b_0/shift_1b_0/n37 ), .ZN(\shifter_0/data_2 [5]) );
  AOI22_X1 \shifter_0/shift_3b_0/shift_1b_0/U39  ( .A1(
        \shifter_0/shift_3b_0/shift_1b_0/n65 ), .A2(\shifter_0/shift_3b_0/n6 ), 
        .B1(\shifter_0/shift_3b_0/n7 ), .B2(
        \shifter_0/shift_3b_0/shift_1b_0/n67 ), .ZN(
        \shifter_0/shift_3b_0/shift_1b_0/n33 ) );
  INV_X1 \shifter_0/shift_3b_0/shift_1b_0/U38  ( .A(
        \shifter_0/shift_3b_0/shift_1b_0/n33 ), .ZN(\shifter_0/data_2 [9]) );
  AOI22_X1 \shifter_0/shift_3b_0/shift_1b_0/U37  ( .A1(
        \shifter_0/shift_3b_0/shift_1b_0/n66 ), .A2(\shifter_0/shift_3b_0/n18 ), .B1(\shifter_0/shift_3b_0/shift_1b_0/n64 ), .B2(\shifter_0/shift_3b_0/n19 ), 
        .ZN(\shifter_0/shift_3b_0/shift_1b_0/n46 ) );
  INV_X1 \shifter_0/shift_3b_0/shift_1b_0/U36  ( .A(
        \shifter_0/shift_3b_0/shift_1b_0/n46 ), .ZN(\shifter_0/data_2 [26]) );
  AOI22_X1 \shifter_0/shift_3b_0/shift_1b_0/U35  ( .A1(
        \shifter_0/shift_3b_0/shift_1b_0/n66 ), .A2(\shifter_0/shift_3b_0/n3 ), 
        .B1(\shifter_0/shift_3b_0/shift_1b_0/n64 ), .B2(
        \shifter_0/shift_3b_0/n18 ), .ZN(\shifter_0/shift_3b_0/shift_1b_0/n45 ) );
  INV_X1 \shifter_0/shift_3b_0/shift_1b_0/U34  ( .A(
        \shifter_0/shift_3b_0/shift_1b_0/n45 ), .ZN(\shifter_0/data_2 [27]) );
  BUF_X1 \shifter_0/shift_3b_0/shift_1b_0/U33  ( .A(
        \shifter_0/shift_3b_0/shift_1b_0/n64 ), .Z(
        \shifter_0/shift_3b_0/shift_1b_0/n67 ) );
  AOI22_X1 \shifter_0/shift_3b_0/shift_1b_0/U32  ( .A1(
        \shifter_0/shift_3b_0/shift_1b_0/n65 ), .A2(\shifter_0/shift_3b_0/n5 ), 
        .B1(\shifter_0/shift_3b_0/shift_1b_0/n64 ), .B2(
        \shifter_0/shift_3b_0/n4 ), .ZN(\shifter_0/shift_3b_0/shift_1b_0/n43 )
         );
  INV_X1 \shifter_0/shift_3b_0/shift_1b_0/U31  ( .A(
        \shifter_0/shift_3b_0/shift_1b_0/n43 ), .ZN(\shifter_0/data_2 [29]) );
  AOI22_X1 \shifter_0/shift_3b_0/shift_1b_0/U30  ( .A1(
        \shifter_0/shift_3b_0/shift_1b_0/n65 ), .A2(\shifter_0/shift_3b_0/n4 ), 
        .B1(\shifter_0/shift_3b_0/shift_1b_0/n64 ), .B2(
        \shifter_0/shift_3b_0/n3 ), .ZN(\shifter_0/shift_3b_0/shift_1b_0/n44 )
         );
  INV_X1 \shifter_0/shift_3b_0/shift_1b_0/U29  ( .A(
        \shifter_0/shift_3b_0/shift_1b_0/n44 ), .ZN(\shifter_0/data_2 [28]) );
  INV_X1 \shifter_0/shift_3b_0/shift_1b_0/U28  ( .A(
        \shifter_0/shift_3b_0/shift_1b_0/n40 ), .ZN(\shifter_0/data_2 [31]) );
  AOI22_X1 \shifter_0/shift_3b_0/shift_1b_0/U27  ( .A1(
        \shifter_0/shift_3b_0/shift_1b_0/n65 ), .A2(\shifter_0/shift_3b_0/n7 ), 
        .B1(\shifter_0/shift_3b_0/shift_1b_0/n64 ), .B2(
        \shifter_0/shift_3b_0/n8 ), .ZN(\shifter_0/shift_3b_0/shift_1b_0/n34 )
         );
  INV_X1 \shifter_0/shift_3b_0/shift_1b_0/U26  ( .A(
        \shifter_0/shift_3b_0/shift_1b_0/n34 ), .ZN(\shifter_0/data_2 [8]) );
  AOI22_X1 \shifter_0/shift_3b_0/shift_1b_0/U25  ( .A1(
        \shifter_0/shift_3b_0/shift_1b_0/n66 ), .A2(\shifter_0/shift_3b_0/n20 ), .B1(\shifter_0/shift_3b_0/shift_1b_0/n64 ), .B2(\shifter_0/shift_3b_0/n21 ), 
        .ZN(\shifter_0/shift_3b_0/shift_1b_0/n48 ) );
  INV_X1 \shifter_0/shift_3b_0/shift_1b_0/U24  ( .A(
        \shifter_0/shift_3b_0/shift_1b_0/n48 ), .ZN(\shifter_0/data_2 [24]) );
  AOI22_X1 \shifter_0/shift_3b_0/shift_1b_0/U23  ( .A1(
        \shifter_0/shift_3b_0/shift_1b_0/n66 ), .A2(\shifter_0/shift_3b_0/n22 ), .B1(\shifter_0/shift_3b_0/shift1 ), .B2(\shifter_0/shift_3b_0/n23 ), .ZN(
        \shifter_0/shift_3b_0/shift_1b_0/n50 ) );
  INV_X1 \shifter_0/shift_3b_0/shift_1b_0/U22  ( .A(
        \shifter_0/shift_3b_0/shift_1b_0/n50 ), .ZN(\shifter_0/data_2 [22]) );
  AOI22_X1 \shifter_0/shift_3b_0/shift_1b_0/U21  ( .A1(
        \shifter_0/shift_3b_0/shift_1b_0/n66 ), .A2(\shifter_0/shift_3b_0/n21 ), .B1(\shifter_0/shift_3b_0/shift1 ), .B2(\shifter_0/shift_3b_0/n22 ), .ZN(
        \shifter_0/shift_3b_0/shift_1b_0/n49 ) );
  INV_X1 \shifter_0/shift_3b_0/shift_1b_0/U20  ( .A(
        \shifter_0/shift_3b_0/shift_1b_0/n49 ), .ZN(\shifter_0/data_2 [23]) );
  AOI22_X1 \shifter_0/shift_3b_0/shift_1b_0/U19  ( .A1(
        \shifter_0/shift_3b_0/shift_1b_0/n66 ), .A2(\shifter_0/shift_3b_0/n25 ), .B1(\shifter_0/shift_3b_0/shift_1b_0/n67 ), .B2(\shifter_0/shift_3b_0/n26 ), 
        .ZN(\shifter_0/shift_3b_0/shift_1b_0/n54 ) );
  INV_X1 \shifter_0/shift_3b_0/shift_1b_0/U18  ( .A(
        \shifter_0/shift_3b_0/shift_1b_0/n54 ), .ZN(\shifter_0/data_2 [19]) );
  AOI22_X1 \shifter_0/shift_3b_0/shift_1b_0/U17  ( .A1(
        \shifter_0/shift_3b_0/shift_1b_0/n66 ), .A2(\shifter_0/shift_3b_0/n24 ), .B1(\shifter_0/shift_3b_0/shift_1b_0/n67 ), .B2(\shifter_0/shift_3b_0/n25 ), 
        .ZN(\shifter_0/shift_3b_0/shift_1b_0/n52 ) );
  INV_X1 \shifter_0/shift_3b_0/shift_1b_0/U16  ( .A(
        \shifter_0/shift_3b_0/shift_1b_0/n52 ), .ZN(\shifter_0/data_2 [20]) );
  AOI22_X1 \shifter_0/shift_3b_0/shift_1b_0/U15  ( .A1(
        \shifter_0/shift_3b_0/shift_1b_0/n66 ), .A2(\shifter_0/shift_3b_0/n23 ), .B1(\shifter_0/shift_3b_0/shift_1b_0/n67 ), .B2(\shifter_0/shift_3b_0/n24 ), 
        .ZN(\shifter_0/shift_3b_0/shift_1b_0/n51 ) );
  INV_X1 \shifter_0/shift_3b_0/shift_1b_0/U14  ( .A(
        \shifter_0/shift_3b_0/shift_1b_0/n51 ), .ZN(\shifter_0/data_2 [21]) );
  AOI22_X1 \shifter_0/shift_3b_0/shift_1b_0/U13  ( .A1(
        \shifter_0/shift_3b_0/shift_1b_0/n65 ), .A2(\shifter_0/shift_3b_0/n29 ), .B1(\shifter_0/shift_3b_0/shift1 ), .B2(\shifter_0/shift_3b_0/n30 ), .ZN(
        \shifter_0/shift_3b_0/shift_1b_0/n58 ) );
  INV_X1 \shifter_0/shift_3b_0/shift_1b_0/U12  ( .A(
        \shifter_0/shift_3b_0/shift_1b_0/n58 ), .ZN(\shifter_0/data_2 [15]) );
  AOI22_X1 \shifter_0/shift_3b_0/shift_1b_0/U11  ( .A1(
        \shifter_0/shift_3b_0/shift_1b_0/n66 ), .A2(\shifter_0/shift_3b_0/n28 ), .B1(\shifter_0/shift_3b_0/shift1 ), .B2(\shifter_0/shift_3b_0/n29 ), .ZN(
        \shifter_0/shift_3b_0/shift_1b_0/n57 ) );
  INV_X1 \shifter_0/shift_3b_0/shift_1b_0/U10  ( .A(
        \shifter_0/shift_3b_0/shift_1b_0/n57 ), .ZN(\shifter_0/data_2 [16]) );
  AOI22_X1 \shifter_0/shift_3b_0/shift_1b_0/U9  ( .A1(
        \shifter_0/shift_3b_0/shift_1b_0/n66 ), .A2(\shifter_0/shift_3b_0/n27 ), .B1(\shifter_0/shift_3b_0/shift1 ), .B2(\shifter_0/shift_3b_0/n28 ), .ZN(
        \shifter_0/shift_3b_0/shift_1b_0/n56 ) );
  INV_X1 \shifter_0/shift_3b_0/shift_1b_0/U8  ( .A(
        \shifter_0/shift_3b_0/shift_1b_0/n56 ), .ZN(\shifter_0/data_2 [17]) );
  AOI22_X1 \shifter_0/shift_3b_0/shift_1b_0/U7  ( .A1(
        \shifter_0/shift_3b_0/shift_1b_0/n66 ), .A2(\shifter_0/shift_3b_0/n26 ), .B1(\shifter_0/shift_3b_0/shift_1b_0/n67 ), .B2(\shifter_0/shift_3b_0/n27 ), 
        .ZN(\shifter_0/shift_3b_0/shift_1b_0/n55 ) );
  INV_X1 \shifter_0/shift_3b_0/shift_1b_0/U6  ( .A(
        \shifter_0/shift_3b_0/shift_1b_0/n55 ), .ZN(\shifter_0/data_2 [18]) );
  AOI22_X1 \shifter_0/shift_3b_0/shift_1b_0/U5  ( .A1(
        \shifter_0/shift_3b_0/shift_1b_0/n66 ), .A2(\shifter_0/shift_3b_0/n19 ), .B1(\shifter_0/shift_3b_0/shift1 ), .B2(\shifter_0/shift_3b_0/n20 ), .ZN(
        \shifter_0/shift_3b_0/shift_1b_0/n47 ) );
  INV_X1 \shifter_0/shift_3b_0/shift_1b_0/U4  ( .A(
        \shifter_0/shift_3b_0/shift_1b_0/n47 ), .ZN(\shifter_0/data_2 [25]) );
  INV_X1 \shifter_0/shift_3b_0/shift_1b_0/U3  ( .A(
        \shifter_0/shift_3b_0/shift1 ), .ZN(
        \shifter_0/shift_3b_0/shift_1b_0/n65 ) );
  INV_X1 \shifter_0/shift_3b_0/shift_1b_0/U2  ( .A(
        \shifter_0/shift_3b_0/shift_1b_0/n64 ), .ZN(
        \shifter_0/shift_3b_0/shift_1b_0/n66 ) );
  INV_X1 \shifter_0/shift_3b_1/U72  ( .A(\shifter_0/n32 ), .ZN(
        \shifter_0/shift_3b_1/n72 ) );
  OAI21_X1 \shifter_0/shift_3b_1/U71  ( .B1(1'b0), .B2(
        \shifter_0/shift_3b_1/n72 ), .A(\shifter_0/shift_3b_1/n35 ), .ZN(
        \shifter_0/shift_3b_1/n61 ) );
  OAI21_X1 \shifter_0/shift_3b_1/U70  ( .B1(\shifter_0/shift_3b_1/n36 ), .B2(
        \shifter_0/shift_3b_1/n72 ), .A(\shifter_0/shift_3b_1/n61 ), .ZN(
        \shifter_0/shift_3b_1/shift1 ) );
  AOI22_X1 \shifter_0/shift_3b_1/U69  ( .A1(\shifter_0/shift_3b_1/n38 ), .A2(
        \shifter_0/data_2 [30]), .B1(\shifter_0/shift_3b_1/n36 ), .B2(
        \shifter_0/data_2 [28]), .ZN(\shifter_0/shift_3b_1/n64 ) );
  INV_X1 \shifter_0/shift_3b_1/U68  ( .A(\shifter_0/shift_3b_1/n64 ), .ZN(
        \shifter_0/shift_3b_1/n4 ) );
  INV_X1 \shifter_0/shift_3b_1/U67  ( .A(\shifter_0/n24 ), .ZN(
        \shifter_0/shift_3b_1/n38 ) );
  INV_X1 \shifter_0/shift_3b_1/U66  ( .A(\shifter_0/data_2 [0]), .ZN(
        \shifter_0/shift_3b_1/n71 ) );
  INV_X1 \shifter_0/shift_3b_1/U65  ( .A(\shifter_0/data_2 [11]), .ZN(
        \shifter_0/shift_3b_1/n69 ) );
  INV_X1 \shifter_0/shift_3b_1/U64  ( .A(\shifter_0/data_2 [10]), .ZN(
        \shifter_0/shift_3b_1/n70 ) );
  INV_X1 \shifter_0/shift_3b_1/U63  ( .A(\shifter_0/data_2 [1]), .ZN(
        \shifter_0/shift_3b_1/n55 ) );
  INV_X1 \shifter_0/shift_3b_1/U62  ( .A(\shifter_0/data_2 [3]), .ZN(
        \shifter_0/shift_3b_1/n45 ) );
  INV_X1 \shifter_0/shift_3b_1/U61  ( .A(\shifter_0/data_2 [4]), .ZN(
        \shifter_0/shift_3b_1/n44 ) );
  INV_X1 \shifter_0/shift_3b_1/U60  ( .A(\shifter_0/data_2 [2]), .ZN(
        \shifter_0/shift_3b_1/n46 ) );
  INV_X1 \shifter_0/shift_3b_1/U59  ( .A(\shifter_0/data_2 [14]), .ZN(
        \shifter_0/shift_3b_1/n66 ) );
  INV_X1 \shifter_0/shift_3b_1/U58  ( .A(\shifter_0/data_2 [13]), .ZN(
        \shifter_0/shift_3b_1/n67 ) );
  INV_X1 \shifter_0/shift_3b_1/U57  ( .A(\shifter_0/data_2 [12]), .ZN(
        \shifter_0/shift_3b_1/n68 ) );
  INV_X1 \shifter_0/shift_3b_1/U56  ( .A(\shifter_0/data_2 [7]), .ZN(
        \shifter_0/shift_3b_1/n41 ) );
  INV_X1 \shifter_0/shift_3b_1/U55  ( .A(\shifter_0/data_2 [6]), .ZN(
        \shifter_0/shift_3b_1/n42 ) );
  INV_X1 \shifter_0/shift_3b_1/U54  ( .A(\shifter_0/data_2 [5]), .ZN(
        \shifter_0/shift_3b_1/n43 ) );
  INV_X1 \shifter_0/shift_3b_1/U53  ( .A(\shifter_0/data_2 [9]), .ZN(
        \shifter_0/shift_3b_1/n39 ) );
  AOI22_X1 \shifter_0/shift_3b_1/U52  ( .A1(\shifter_0/shift_3b_1/n38 ), .A2(
        \shifter_0/data_2 [31]), .B1(\shifter_0/shift_3b_1/n36 ), .B2(
        \shifter_0/data_2 [29]), .ZN(\shifter_0/shift_3b_1/n65 ) );
  INV_X1 \shifter_0/shift_3b_1/U51  ( .A(\shifter_0/shift_3b_1/n65 ), .ZN(
        \shifter_0/shift_3b_1/n14 ) );
  INV_X1 \shifter_0/shift_3b_1/U50  ( .A(\shifter_0/data_2 [8]), .ZN(
        \shifter_0/shift_3b_1/n40 ) );
  INV_X1 \shifter_0/shift_3b_1/U49  ( .A(\shifter_0/data_2 [24]), .ZN(
        \shifter_0/shift_3b_1/n50 ) );
  INV_X1 \shifter_0/shift_3b_1/U48  ( .A(\shifter_0/data_2 [22]), .ZN(
        \shifter_0/shift_3b_1/n52 ) );
  INV_X1 \shifter_0/shift_3b_1/U47  ( .A(\shifter_0/data_2 [23]), .ZN(
        \shifter_0/shift_3b_1/n51 ) );
  INV_X1 \shifter_0/shift_3b_1/U46  ( .A(\shifter_0/data_2 [19]), .ZN(
        \shifter_0/shift_3b_1/n56 ) );
  INV_X1 \shifter_0/shift_3b_1/U45  ( .A(\shifter_0/data_2 [20]), .ZN(
        \shifter_0/shift_3b_1/n54 ) );
  INV_X1 \shifter_0/shift_3b_1/U44  ( .A(\shifter_0/data_2 [21]), .ZN(
        \shifter_0/shift_3b_1/n53 ) );
  INV_X1 \shifter_0/shift_3b_1/U43  ( .A(\shifter_0/data_2 [15]), .ZN(
        \shifter_0/shift_3b_1/n60 ) );
  INV_X1 \shifter_0/shift_3b_1/U42  ( .A(\shifter_0/data_2 [16]), .ZN(
        \shifter_0/shift_3b_1/n59 ) );
  INV_X1 \shifter_0/shift_3b_1/U41  ( .A(\shifter_0/data_2 [17]), .ZN(
        \shifter_0/shift_3b_1/n58 ) );
  INV_X1 \shifter_0/shift_3b_1/U40  ( .A(\shifter_0/data_2 [18]), .ZN(
        \shifter_0/shift_3b_1/n57 ) );
  INV_X1 \shifter_0/shift_3b_1/U39  ( .A(\shifter_0/data_2 [25]), .ZN(
        \shifter_0/shift_3b_1/n49 ) );
  AOI22_X1 \shifter_0/shift_3b_1/U38  ( .A1(\shifter_0/shift_3b_1/n38 ), .A2(
        \shifter_0/data_2 [28]), .B1(\shifter_0/shift_3b_1/n36 ), .B2(
        \shifter_0/data_2 [26]), .ZN(\shifter_0/shift_3b_1/n62 ) );
  INV_X1 \shifter_0/shift_3b_1/U37  ( .A(\shifter_0/shift_3b_1/n62 ), .ZN(
        \shifter_0/shift_3b_1/n2 ) );
  AOI22_X1 \shifter_0/shift_3b_1/U36  ( .A1(\shifter_0/shift_3b_1/n38 ), .A2(
        \shifter_0/data_2 [29]), .B1(\shifter_0/shift_3b_1/n36 ), .B2(
        \shifter_0/data_2 [27]), .ZN(\shifter_0/shift_3b_1/n63 ) );
  INV_X1 \shifter_0/shift_3b_1/U35  ( .A(\shifter_0/shift_3b_1/n63 ), .ZN(
        \shifter_0/shift_3b_1/n3 ) );
  NOR2_X1 \shifter_0/shift_3b_1/U34  ( .A1(\shifter_0/shift_3b_1/n35 ), .A2(
        \shifter_0/shift_3b_1/n71 ), .ZN(\shifter_0/shift_3b_1/data1 [0]) );
  NOR2_X1 \shifter_0/shift_3b_1/U33  ( .A1(\shifter_0/shift_3b_1/n35 ), .A2(
        \shifter_0/shift_3b_1/n55 ), .ZN(\shifter_0/shift_3b_1/data1 [1]) );
  OAI22_X1 \shifter_0/shift_3b_1/U32  ( .A1(\shifter_0/shift_3b_1/n35 ), .A2(
        \shifter_0/shift_3b_1/n40 ), .B1(\shifter_0/shift_3b_1/n38 ), .B2(
        \shifter_0/shift_3b_1/n42 ), .ZN(\shifter_0/shift_3b_1/n8 ) );
  OAI22_X1 \shifter_0/shift_3b_1/U31  ( .A1(\shifter_0/shift_3b_1/n36 ), .A2(
        \shifter_0/shift_3b_1/n54 ), .B1(\shifter_0/shift_3b_1/n38 ), .B2(
        \shifter_0/shift_3b_1/n57 ), .ZN(\shifter_0/shift_3b_1/n26 ) );
  OAI22_X1 \shifter_0/shift_3b_1/U30  ( .A1(\shifter_0/shift_3b_1/n36 ), .A2(
        \shifter_0/shift_3b_1/n50 ), .B1(\shifter_0/shift_3b_1/n38 ), .B2(
        \shifter_0/shift_3b_1/n52 ), .ZN(\shifter_0/shift_3b_1/n22 ) );
  OAI22_X1 \shifter_0/shift_3b_1/U29  ( .A1(\shifter_0/shift_3b_1/n36 ), .A2(
        \shifter_0/shift_3b_1/n53 ), .B1(\shifter_0/shift_3b_1/n38 ), .B2(
        \shifter_0/shift_3b_1/n56 ), .ZN(\shifter_0/shift_3b_1/n25 ) );
  OAI22_X1 \shifter_0/shift_3b_1/U28  ( .A1(\shifter_0/shift_3b_1/n36 ), .A2(
        \shifter_0/shift_3b_1/n52 ), .B1(\shifter_0/shift_3b_1/n38 ), .B2(
        \shifter_0/shift_3b_1/n54 ), .ZN(\shifter_0/shift_3b_1/n24 ) );
  OAI22_X1 \shifter_0/shift_3b_1/U27  ( .A1(\shifter_0/shift_3b_1/n36 ), .A2(
        \shifter_0/shift_3b_1/n51 ), .B1(\shifter_0/shift_3b_1/n38 ), .B2(
        \shifter_0/shift_3b_1/n53 ), .ZN(\shifter_0/shift_3b_1/n23 ) );
  OAI22_X1 \shifter_0/shift_3b_1/U26  ( .A1(\shifter_0/shift_3b_1/n36 ), .A2(
        \shifter_0/shift_3b_1/n56 ), .B1(\shifter_0/shift_3b_1/n38 ), .B2(
        \shifter_0/shift_3b_1/n58 ), .ZN(\shifter_0/shift_3b_1/n27 ) );
  OAI22_X1 \shifter_0/shift_3b_1/U25  ( .A1(\shifter_0/shift_3b_1/n36 ), .A2(
        \shifter_0/shift_3b_1/n67 ), .B1(\shifter_0/shift_3b_1/n38 ), .B2(
        \shifter_0/shift_3b_1/n69 ), .ZN(\shifter_0/shift_3b_1/n33 ) );
  OAI22_X1 \shifter_0/shift_3b_1/U24  ( .A1(\shifter_0/shift_3b_1/n36 ), .A2(
        \shifter_0/shift_3b_1/n59 ), .B1(\shifter_0/shift_3b_1/n37 ), .B2(
        \shifter_0/shift_3b_1/n66 ), .ZN(\shifter_0/shift_3b_1/n30 ) );
  OAI22_X1 \shifter_0/shift_3b_1/U23  ( .A1(\shifter_0/shift_3b_1/n35 ), .A2(
        \shifter_0/shift_3b_1/n60 ), .B1(\shifter_0/shift_3b_1/n37 ), .B2(
        \shifter_0/shift_3b_1/n67 ), .ZN(\shifter_0/shift_3b_1/n31 ) );
  OAI22_X1 \shifter_0/shift_3b_1/U22  ( .A1(\shifter_0/shift_3b_1/n35 ), .A2(
        \shifter_0/shift_3b_1/n66 ), .B1(\shifter_0/shift_3b_1/n37 ), .B2(
        \shifter_0/shift_3b_1/n68 ), .ZN(\shifter_0/shift_3b_1/n32 ) );
  OAI22_X1 \shifter_0/shift_3b_1/U21  ( .A1(\shifter_0/shift_3b_1/n36 ), .A2(
        \shifter_0/shift_3b_1/n58 ), .B1(\shifter_0/shift_3b_1/n38 ), .B2(
        \shifter_0/shift_3b_1/n60 ), .ZN(\shifter_0/shift_3b_1/n29 ) );
  OAI22_X1 \shifter_0/shift_3b_1/U20  ( .A1(\shifter_0/shift_3b_1/n36 ), .A2(
        \shifter_0/shift_3b_1/n57 ), .B1(\shifter_0/shift_3b_1/n38 ), .B2(
        \shifter_0/shift_3b_1/n59 ), .ZN(\shifter_0/shift_3b_1/n28 ) );
  OAI22_X1 \shifter_0/shift_3b_1/U19  ( .A1(\shifter_0/shift_3b_1/n35 ), .A2(
        \shifter_0/shift_3b_1/n68 ), .B1(\shifter_0/shift_3b_1/n38 ), .B2(
        \shifter_0/shift_3b_1/n70 ), .ZN(\shifter_0/shift_3b_1/n34 ) );
  INV_X1 \shifter_0/shift_3b_1/U18  ( .A(\shifter_0/data_2 [26]), .ZN(
        \shifter_0/shift_3b_1/n48 ) );
  OAI22_X1 \shifter_0/shift_3b_1/U17  ( .A1(\shifter_0/shift_3b_1/n36 ), .A2(
        \shifter_0/shift_3b_1/n48 ), .B1(\shifter_0/shift_3b_1/n38 ), .B2(
        \shifter_0/shift_3b_1/n50 ), .ZN(\shifter_0/shift_3b_1/n20 ) );
  OAI22_X1 \shifter_0/shift_3b_1/U16  ( .A1(\shifter_0/shift_3b_1/n36 ), .A2(
        \shifter_0/shift_3b_1/n49 ), .B1(\shifter_0/shift_3b_1/n38 ), .B2(
        \shifter_0/shift_3b_1/n51 ), .ZN(\shifter_0/shift_3b_1/n21 ) );
  OAI22_X1 \shifter_0/shift_3b_1/U15  ( .A1(\shifter_0/shift_3b_1/n35 ), .A2(
        \shifter_0/shift_3b_1/n41 ), .B1(\shifter_0/shift_3b_1/n38 ), .B2(
        \shifter_0/shift_3b_1/n43 ), .ZN(\shifter_0/shift_3b_1/n9 ) );
  OAI22_X1 \shifter_0/shift_3b_1/U14  ( .A1(\shifter_0/shift_3b_1/n36 ), .A2(
        \shifter_0/shift_3b_1/n43 ), .B1(\shifter_0/shift_3b_1/n38 ), .B2(
        \shifter_0/shift_3b_1/n45 ), .ZN(\shifter_0/shift_3b_1/n11 ) );
  OAI22_X1 \shifter_0/shift_3b_1/U13  ( .A1(\shifter_0/shift_3b_1/n35 ), .A2(
        \shifter_0/shift_3b_1/n42 ), .B1(\shifter_0/shift_3b_1/n38 ), .B2(
        \shifter_0/shift_3b_1/n44 ), .ZN(\shifter_0/shift_3b_1/n10 ) );
  OAI22_X1 \shifter_0/shift_3b_1/U12  ( .A1(\shifter_0/n24 ), .A2(
        \shifter_0/shift_3b_1/n46 ), .B1(\shifter_0/shift_3b_1/n38 ), .B2(
        \shifter_0/shift_3b_1/n71 ), .ZN(\shifter_0/shift_3b_1/n16 ) );
  OAI22_X1 \shifter_0/shift_3b_1/U11  ( .A1(\shifter_0/shift_3b_1/n36 ), .A2(
        \shifter_0/shift_3b_1/n44 ), .B1(\shifter_0/shift_3b_1/n38 ), .B2(
        \shifter_0/shift_3b_1/n46 ), .ZN(\shifter_0/shift_3b_1/n12 ) );
  OAI22_X1 \shifter_0/shift_3b_1/U10  ( .A1(\shifter_0/shift_3b_1/n36 ), .A2(
        \shifter_0/shift_3b_1/n45 ), .B1(\shifter_0/shift_3b_1/n38 ), .B2(
        \shifter_0/shift_3b_1/n55 ), .ZN(\shifter_0/shift_3b_1/n13 ) );
  INV_X1 \shifter_0/shift_3b_1/U9  ( .A(\shifter_0/data_2 [27]), .ZN(
        \shifter_0/shift_3b_1/n47 ) );
  OAI22_X1 \shifter_0/shift_3b_1/U8  ( .A1(\shifter_0/n24 ), .A2(
        \shifter_0/shift_3b_1/n47 ), .B1(\shifter_0/shift_3b_1/n38 ), .B2(
        \shifter_0/shift_3b_1/n49 ), .ZN(\shifter_0/shift_3b_1/n19 ) );
  OAI22_X1 \shifter_0/shift_3b_1/U7  ( .A1(\shifter_0/shift_3b_1/n37 ), .A2(
        \shifter_0/shift_3b_1/n40 ), .B1(\shifter_0/shift_3b_1/n35 ), .B2(
        \shifter_0/shift_3b_1/n70 ), .ZN(\shifter_0/shift_3b_1/n7 ) );
  OAI22_X1 \shifter_0/shift_3b_1/U6  ( .A1(\shifter_0/shift_3b_1/n35 ), .A2(
        \shifter_0/shift_3b_1/n39 ), .B1(\shifter_0/shift_3b_1/n38 ), .B2(
        \shifter_0/shift_3b_1/n41 ), .ZN(\shifter_0/shift_3b_1/n6 ) );
  OAI22_X1 \shifter_0/shift_3b_1/U5  ( .A1(\shifter_0/shift_3b_1/n37 ), .A2(
        \shifter_0/shift_3b_1/n39 ), .B1(\shifter_0/shift_3b_1/n35 ), .B2(
        \shifter_0/shift_3b_1/n69 ), .ZN(\shifter_0/shift_3b_1/n5 ) );
  INV_X1 \shifter_0/shift_3b_1/U4  ( .A(\shifter_0/shift_3b_1/n37 ), .ZN(
        \shifter_0/shift_3b_1/n36 ) );
  INV_X1 \shifter_0/shift_3b_1/U3  ( .A(\shifter_0/shift_3b_1/n37 ), .ZN(
        \shifter_0/shift_3b_1/n35 ) );
  CLKBUF_X1 \shifter_0/shift_3b_1/U2  ( .A(\shifter_0/shift_3b_1/n38 ), .Z(
        \shifter_0/shift_3b_1/n37 ) );
  BUF_X1 \shifter_0/shift_3b_1/shift_1b_0/U69  ( .A(
        \shifter_0/shift_3b_1/shift1 ), .Z(
        \shifter_0/shift_3b_1/shift_1b_0/n64 ) );
  AOI22_X1 \shifter_0/shift_3b_1/shift_1b_0/U68  ( .A1(
        \shifter_0/shift_3b_1/shift_1b_0/n65 ), .A2(\shifter_0/shift_3b_1/n4 ), 
        .B1(\shifter_0/shift_3b_1/shift_1b_0/n64 ), .B2(
        \shifter_0/shift_3b_1/n3 ), .ZN(\shifter_0/shift_3b_1/shift_1b_0/n91 )
         );
  INV_X1 \shifter_0/shift_3b_1/shift_1b_0/U67  ( .A(
        \shifter_0/shift_3b_1/shift_1b_0/n91 ), .ZN(\shifter_0/data_3 [30]) );
  BUF_X1 \shifter_0/shift_3b_1/shift_1b_0/U66  ( .A(
        \shifter_0/shift_3b_1/shift_1b_0/n64 ), .Z(
        \shifter_0/shift_3b_1/shift_1b_0/n67 ) );
  AOI22_X1 \shifter_0/shift_3b_1/shift_1b_0/U65  ( .A1(
        \shifter_0/shift_3b_1/shift_1b_0/n65 ), .A2(\shifter_0/shift_3b_1/n14 ), .B1(\shifter_0/shift_3b_1/shift_1b_0/n64 ), .B2(\shifter_0/shift_3b_1/n4 ), 
        .ZN(\shifter_0/shift_3b_1/shift_1b_0/n92 ) );
  AOI22_X1 \shifter_0/shift_3b_1/shift_1b_0/U64  ( .A1(
        \shifter_0/shift_3b_1/shift_1b_0/n65 ), .A2(\shifter_0/shift_3b_1/n6 ), 
        .B1(\shifter_0/shift_3b_1/n8 ), .B2(
        \shifter_0/shift_3b_1/shift_1b_0/n68 ), .ZN(
        \shifter_0/shift_3b_1/shift_1b_0/n99 ) );
  INV_X1 \shifter_0/shift_3b_1/shift_1b_0/U63  ( .A(
        \shifter_0/shift_3b_1/shift_1b_0/n99 ), .ZN(\shifter_0/data_3 [9]) );
  INV_X1 \shifter_0/shift_3b_1/shift_1b_0/U62  ( .A(
        \shifter_0/shift_3b_1/shift_1b_0/n92 ), .ZN(\shifter_0/data_3 [31]) );
  AOI22_X1 \shifter_0/shift_3b_1/shift_1b_0/U61  ( .A1(
        \shifter_0/shift_3b_1/shift_1b_0/n65 ), .A2(\shifter_0/shift_3b_1/n5 ), 
        .B1(\shifter_0/shift_3b_1/shift_1b_0/n68 ), .B2(
        \shifter_0/shift_3b_1/n7 ), .ZN(\shifter_0/shift_3b_1/shift_1b_0/n70 )
         );
  INV_X1 \shifter_0/shift_3b_1/shift_1b_0/U60  ( .A(
        \shifter_0/shift_3b_1/shift_1b_0/n70 ), .ZN(\shifter_0/data_3 [11]) );
  AOI22_X1 \shifter_0/shift_3b_1/shift_1b_0/U59  ( .A1(
        \shifter_0/shift_3b_1/shift_1b_0/n65 ), .A2(\shifter_0/shift_3b_1/n34 ), .B1(\shifter_0/shift_3b_1/shift_1b_0/n68 ), .B2(\shifter_0/shift_3b_1/n5 ), 
        .ZN(\shifter_0/shift_3b_1/shift_1b_0/n71 ) );
  INV_X1 \shifter_0/shift_3b_1/shift_1b_0/U58  ( .A(
        \shifter_0/shift_3b_1/shift_1b_0/n71 ), .ZN(\shifter_0/data_3 [12]) );
  AOI22_X1 \shifter_0/shift_3b_1/shift_1b_0/U57  ( .A1(
        \shifter_0/shift_3b_1/shift_1b_0/n65 ), .A2(\shifter_0/shift_3b_1/n33 ), .B1(\shifter_0/shift_3b_1/shift_1b_0/n68 ), .B2(\shifter_0/shift_3b_1/n34 ), 
        .ZN(\shifter_0/shift_3b_1/shift_1b_0/n72 ) );
  INV_X1 \shifter_0/shift_3b_1/shift_1b_0/U56  ( .A(
        \shifter_0/shift_3b_1/shift_1b_0/n72 ), .ZN(\shifter_0/data_3 [13]) );
  AOI22_X1 \shifter_0/shift_3b_1/shift_1b_0/U55  ( .A1(
        \shifter_0/shift_3b_1/shift_1b_0/n64 ), .A2(\shifter_0/shift_3b_1/n6 ), 
        .B1(\shifter_0/shift_3b_1/shift_1b_0/n66 ), .B2(
        \shifter_0/shift_3b_1/n7 ), .ZN(\shifter_0/shift_3b_1/shift_1b_0/n69 )
         );
  INV_X1 \shifter_0/shift_3b_1/shift_1b_0/U54  ( .A(
        \shifter_0/shift_3b_1/shift_1b_0/n69 ), .ZN(\shifter_0/data_3 [10]) );
  AOI22_X1 \shifter_0/shift_3b_1/shift_1b_0/U53  ( .A1(
        \shifter_0/shift_3b_1/shift_1b_0/n65 ), .A2(\shifter_0/shift_3b_1/n8 ), 
        .B1(\shifter_0/shift_3b_1/shift_1b_0/n67 ), .B2(
        \shifter_0/shift_3b_1/n9 ), .ZN(\shifter_0/shift_3b_1/shift_1b_0/n98 )
         );
  INV_X1 \shifter_0/shift_3b_1/shift_1b_0/U52  ( .A(
        \shifter_0/shift_3b_1/shift_1b_0/n98 ), .ZN(\shifter_0/data_3 [8]) );
  AOI22_X1 \shifter_0/shift_3b_1/shift_1b_0/U51  ( .A1(
        \shifter_0/shift_3b_1/shift_1b_0/n66 ), .A2(
        \shifter_0/shift_3b_1/data1 [1]), .B1(
        \shifter_0/shift_3b_1/shift_1b_0/n64 ), .B2(
        \shifter_0/shift_3b_1/data1 [0]), .ZN(
        \shifter_0/shift_3b_1/shift_1b_0/n79 ) );
  INV_X1 \shifter_0/shift_3b_1/shift_1b_0/U50  ( .A(
        \shifter_0/shift_3b_1/shift_1b_0/n79 ), .ZN(\shifter_0/data_3 [1]) );
  AOI22_X1 \shifter_0/shift_3b_1/shift_1b_0/U49  ( .A1(
        \shifter_0/shift_3b_1/shift_1b_0/n65 ), .A2(\shifter_0/shift_3b_1/n9 ), 
        .B1(\shifter_0/shift_3b_1/shift_1b_0/n67 ), .B2(
        \shifter_0/shift_3b_1/n10 ), .ZN(\shifter_0/shift_3b_1/shift_1b_0/n97 ) );
  INV_X1 \shifter_0/shift_3b_1/shift_1b_0/U48  ( .A(
        \shifter_0/shift_3b_1/shift_1b_0/n97 ), .ZN(\shifter_0/data_3 [7]) );
  AOI22_X1 \shifter_0/shift_3b_1/shift_1b_0/U47  ( .A1(
        \shifter_0/shift_3b_1/shift_1b_0/n65 ), .A2(\shifter_0/shift_3b_1/n10 ), .B1(\shifter_0/shift_3b_1/shift_1b_0/n67 ), .B2(\shifter_0/shift_3b_1/n11 ), 
        .ZN(\shifter_0/shift_3b_1/shift_1b_0/n96 ) );
  INV_X1 \shifter_0/shift_3b_1/shift_1b_0/U46  ( .A(
        \shifter_0/shift_3b_1/shift_1b_0/n96 ), .ZN(\shifter_0/data_3 [6]) );
  AOI22_X1 \shifter_0/shift_3b_1/shift_1b_0/U45  ( .A1(
        \shifter_0/shift_3b_1/shift_1b_0/n65 ), .A2(\shifter_0/shift_3b_1/n16 ), .B1(\shifter_0/shift_3b_1/shift_1b_0/n68 ), .B2(
        \shifter_0/shift_3b_1/data1 [1]), .ZN(
        \shifter_0/shift_3b_1/shift_1b_0/n90 ) );
  INV_X1 \shifter_0/shift_3b_1/shift_1b_0/U44  ( .A(
        \shifter_0/shift_3b_1/shift_1b_0/n90 ), .ZN(\shifter_0/data_3 [2]) );
  AOI22_X1 \shifter_0/shift_3b_1/shift_1b_0/U43  ( .A1(
        \shifter_0/shift_3b_1/shift_1b_0/n65 ), .A2(\shifter_0/shift_3b_1/n13 ), .B1(\shifter_0/shift_3b_1/shift_1b_0/n67 ), .B2(\shifter_0/shift_3b_1/n16 ), 
        .ZN(\shifter_0/shift_3b_1/shift_1b_0/n93 ) );
  INV_X1 \shifter_0/shift_3b_1/shift_1b_0/U42  ( .A(
        \shifter_0/shift_3b_1/shift_1b_0/n93 ), .ZN(\shifter_0/data_3 [3]) );
  AOI22_X1 \shifter_0/shift_3b_1/shift_1b_0/U41  ( .A1(
        \shifter_0/shift_3b_1/shift_1b_0/n65 ), .A2(\shifter_0/shift_3b_1/n11 ), .B1(\shifter_0/shift_3b_1/shift_1b_0/n67 ), .B2(\shifter_0/shift_3b_1/n12 ), 
        .ZN(\shifter_0/shift_3b_1/shift_1b_0/n95 ) );
  INV_X1 \shifter_0/shift_3b_1/shift_1b_0/U40  ( .A(
        \shifter_0/shift_3b_1/shift_1b_0/n95 ), .ZN(\shifter_0/data_3 [5]) );
  AOI22_X1 \shifter_0/shift_3b_1/shift_1b_0/U39  ( .A1(
        \shifter_0/shift_3b_1/shift_1b_0/n65 ), .A2(\shifter_0/shift_3b_1/n12 ), .B1(\shifter_0/shift_3b_1/shift_1b_0/n67 ), .B2(\shifter_0/shift_3b_1/n13 ), 
        .ZN(\shifter_0/shift_3b_1/shift_1b_0/n94 ) );
  INV_X1 \shifter_0/shift_3b_1/shift_1b_0/U38  ( .A(
        \shifter_0/shift_3b_1/shift_1b_0/n94 ), .ZN(\shifter_0/data_3 [4]) );
  AOI22_X1 \shifter_0/shift_3b_1/shift_1b_0/U37  ( .A1(
        \shifter_0/shift_3b_1/shift_1b_0/n65 ), .A2(\shifter_0/shift_3b_1/n32 ), .B1(\shifter_0/shift_3b_1/shift_1b_0/n67 ), .B2(\shifter_0/shift_3b_1/n33 ), 
        .ZN(\shifter_0/shift_3b_1/shift_1b_0/n73 ) );
  INV_X1 \shifter_0/shift_3b_1/shift_1b_0/U36  ( .A(
        \shifter_0/shift_3b_1/shift_1b_0/n73 ), .ZN(\shifter_0/data_3 [14]) );
  AOI22_X1 \shifter_0/shift_3b_1/shift_1b_0/U35  ( .A1(
        \shifter_0/shift_3b_1/shift_1b_0/n66 ), .A2(\shifter_0/shift_3b_1/n29 ), .B1(\shifter_0/shift_3b_1/shift_1b_0/n67 ), .B2(\shifter_0/shift_3b_1/n30 ), 
        .ZN(\shifter_0/shift_3b_1/shift_1b_0/n76 ) );
  INV_X1 \shifter_0/shift_3b_1/shift_1b_0/U34  ( .A(
        \shifter_0/shift_3b_1/shift_1b_0/n76 ), .ZN(\shifter_0/data_3 [17]) );
  AOI22_X1 \shifter_0/shift_3b_1/shift_1b_0/U33  ( .A1(
        \shifter_0/shift_3b_1/shift_1b_0/n66 ), .A2(\shifter_0/shift_3b_1/n30 ), .B1(\shifter_0/shift_3b_1/shift_1b_0/n67 ), .B2(\shifter_0/shift_3b_1/n31 ), 
        .ZN(\shifter_0/shift_3b_1/shift_1b_0/n75 ) );
  INV_X1 \shifter_0/shift_3b_1/shift_1b_0/U32  ( .A(
        \shifter_0/shift_3b_1/shift_1b_0/n75 ), .ZN(\shifter_0/data_3 [16]) );
  AOI22_X1 \shifter_0/shift_3b_1/shift_1b_0/U31  ( .A1(
        \shifter_0/shift_3b_1/shift_1b_0/n66 ), .A2(\shifter_0/shift_3b_1/n31 ), .B1(\shifter_0/shift_3b_1/shift_1b_0/n67 ), .B2(\shifter_0/shift_3b_1/n32 ), 
        .ZN(\shifter_0/shift_3b_1/shift_1b_0/n74 ) );
  INV_X1 \shifter_0/shift_3b_1/shift_1b_0/U30  ( .A(
        \shifter_0/shift_3b_1/shift_1b_0/n74 ), .ZN(\shifter_0/data_3 [15]) );
  AOI22_X1 \shifter_0/shift_3b_1/shift_1b_0/U29  ( .A1(
        \shifter_0/shift_3b_1/shift_1b_0/n66 ), .A2(\shifter_0/shift_3b_1/n28 ), .B1(\shifter_0/shift_3b_1/shift_1b_0/n67 ), .B2(\shifter_0/shift_3b_1/n29 ), 
        .ZN(\shifter_0/shift_3b_1/shift_1b_0/n77 ) );
  INV_X1 \shifter_0/shift_3b_1/shift_1b_0/U28  ( .A(
        \shifter_0/shift_3b_1/shift_1b_0/n77 ), .ZN(\shifter_0/data_3 [18]) );
  AOI22_X1 \shifter_0/shift_3b_1/shift_1b_0/U27  ( .A1(
        \shifter_0/shift_3b_1/shift_1b_0/n66 ), .A2(\shifter_0/shift_3b_1/n27 ), .B1(\shifter_0/shift_3b_1/shift_1b_0/n68 ), .B2(\shifter_0/shift_3b_1/n28 ), 
        .ZN(\shifter_0/shift_3b_1/shift_1b_0/n78 ) );
  INV_X1 \shifter_0/shift_3b_1/shift_1b_0/U26  ( .A(
        \shifter_0/shift_3b_1/shift_1b_0/n78 ), .ZN(\shifter_0/data_3 [19]) );
  AOI22_X1 \shifter_0/shift_3b_1/shift_1b_0/U25  ( .A1(
        \shifter_0/shift_3b_1/shift_1b_0/n66 ), .A2(\shifter_0/shift_3b_1/n26 ), .B1(\shifter_0/shift_3b_1/shift_1b_0/n64 ), .B2(\shifter_0/shift_3b_1/n27 ), 
        .ZN(\shifter_0/shift_3b_1/shift_1b_0/n80 ) );
  INV_X1 \shifter_0/shift_3b_1/shift_1b_0/U24  ( .A(
        \shifter_0/shift_3b_1/shift_1b_0/n80 ), .ZN(\shifter_0/data_3 [20]) );
  AOI22_X1 \shifter_0/shift_3b_1/shift_1b_0/U23  ( .A1(
        \shifter_0/shift_3b_1/shift_1b_0/n66 ), .A2(\shifter_0/shift_3b_1/n25 ), .B1(\shifter_0/shift_3b_1/shift_1b_0/n64 ), .B2(\shifter_0/shift_3b_1/n26 ), 
        .ZN(\shifter_0/shift_3b_1/shift_1b_0/n81 ) );
  INV_X1 \shifter_0/shift_3b_1/shift_1b_0/U22  ( .A(
        \shifter_0/shift_3b_1/shift_1b_0/n81 ), .ZN(\shifter_0/data_3 [21]) );
  AOI22_X1 \shifter_0/shift_3b_1/shift_1b_0/U21  ( .A1(
        \shifter_0/shift_3b_1/shift_1b_0/n66 ), .A2(\shifter_0/shift_3b_1/n24 ), .B1(\shifter_0/shift_3b_1/shift_1b_0/n64 ), .B2(\shifter_0/shift_3b_1/n25 ), 
        .ZN(\shifter_0/shift_3b_1/shift_1b_0/n82 ) );
  INV_X1 \shifter_0/shift_3b_1/shift_1b_0/U20  ( .A(
        \shifter_0/shift_3b_1/shift_1b_0/n82 ), .ZN(\shifter_0/data_3 [22]) );
  AOI22_X1 \shifter_0/shift_3b_1/shift_1b_0/U19  ( .A1(
        \shifter_0/shift_3b_1/shift_1b_0/n66 ), .A2(\shifter_0/shift_3b_1/n23 ), .B1(\shifter_0/shift_3b_1/shift_1b_0/n64 ), .B2(\shifter_0/shift_3b_1/n24 ), 
        .ZN(\shifter_0/shift_3b_1/shift_1b_0/n83 ) );
  INV_X1 \shifter_0/shift_3b_1/shift_1b_0/U18  ( .A(
        \shifter_0/shift_3b_1/shift_1b_0/n83 ), .ZN(\shifter_0/data_3 [23]) );
  AOI22_X1 \shifter_0/shift_3b_1/shift_1b_0/U17  ( .A1(
        \shifter_0/shift_3b_1/shift_1b_0/n66 ), .A2(\shifter_0/shift_3b_1/n22 ), .B1(\shifter_0/shift_3b_1/shift_1b_0/n64 ), .B2(\shifter_0/shift_3b_1/n23 ), 
        .ZN(\shifter_0/shift_3b_1/shift_1b_0/n84 ) );
  INV_X1 \shifter_0/shift_3b_1/shift_1b_0/U16  ( .A(
        \shifter_0/shift_3b_1/shift_1b_0/n84 ), .ZN(\shifter_0/data_3 [24]) );
  AOI22_X1 \shifter_0/shift_3b_1/shift_1b_0/U15  ( .A1(
        \shifter_0/shift_3b_1/shift_1b_0/n66 ), .A2(\shifter_0/shift_3b_1/n21 ), .B1(\shifter_0/shift_3b_1/shift_1b_0/n64 ), .B2(\shifter_0/shift_3b_1/n22 ), 
        .ZN(\shifter_0/shift_3b_1/shift_1b_0/n85 ) );
  INV_X1 \shifter_0/shift_3b_1/shift_1b_0/U14  ( .A(
        \shifter_0/shift_3b_1/shift_1b_0/n85 ), .ZN(\shifter_0/data_3 [25]) );
  AOI22_X1 \shifter_0/shift_3b_1/shift_1b_0/U13  ( .A1(
        \shifter_0/shift_3b_1/shift_1b_0/n66 ), .A2(\shifter_0/shift_3b_1/n19 ), .B1(\shifter_0/shift_3b_1/shift_1b_0/n64 ), .B2(\shifter_0/shift_3b_1/n20 ), 
        .ZN(\shifter_0/shift_3b_1/shift_1b_0/n87 ) );
  INV_X1 \shifter_0/shift_3b_1/shift_1b_0/U12  ( .A(
        \shifter_0/shift_3b_1/shift_1b_0/n87 ), .ZN(\shifter_0/data_3 [27]) );
  AOI22_X1 \shifter_0/shift_3b_1/shift_1b_0/U11  ( .A1(
        \shifter_0/shift_3b_1/shift_1b_0/n66 ), .A2(\shifter_0/shift_3b_1/n20 ), .B1(\shifter_0/shift_3b_1/shift_1b_0/n64 ), .B2(\shifter_0/shift_3b_1/n21 ), 
        .ZN(\shifter_0/shift_3b_1/shift_1b_0/n86 ) );
  INV_X1 \shifter_0/shift_3b_1/shift_1b_0/U10  ( .A(
        \shifter_0/shift_3b_1/shift_1b_0/n86 ), .ZN(\shifter_0/data_3 [26]) );
  AOI22_X1 \shifter_0/shift_3b_1/shift_1b_0/U9  ( .A1(
        \shifter_0/shift_3b_1/shift_1b_0/n65 ), .A2(\shifter_0/shift_3b_1/n2 ), 
        .B1(\shifter_0/shift_3b_1/shift_1b_0/n64 ), .B2(
        \shifter_0/shift_3b_1/n19 ), .ZN(\shifter_0/shift_3b_1/shift_1b_0/n88 ) );
  INV_X1 \shifter_0/shift_3b_1/shift_1b_0/U8  ( .A(
        \shifter_0/shift_3b_1/shift_1b_0/n88 ), .ZN(\shifter_0/data_3 [28]) );
  AOI22_X1 \shifter_0/shift_3b_1/shift_1b_0/U7  ( .A1(
        \shifter_0/shift_3b_1/shift_1b_0/n65 ), .A2(\shifter_0/shift_3b_1/n3 ), 
        .B1(\shifter_0/shift_3b_1/shift_1b_0/n64 ), .B2(
        \shifter_0/shift_3b_1/n2 ), .ZN(\shifter_0/shift_3b_1/shift_1b_0/n89 )
         );
  INV_X1 \shifter_0/shift_3b_1/shift_1b_0/U6  ( .A(
        \shifter_0/shift_3b_1/shift_1b_0/n89 ), .ZN(\shifter_0/data_3 [29]) );
  INV_X1 \shifter_0/shift_3b_1/shift_1b_0/U5  ( .A(
        \shifter_0/shift_3b_1/shift1 ), .ZN(
        \shifter_0/shift_3b_1/shift_1b_0/n66 ) );
  INV_X1 \shifter_0/shift_3b_1/shift_1b_0/U4  ( .A(
        \shifter_0/shift_3b_1/shift1 ), .ZN(
        \shifter_0/shift_3b_1/shift_1b_0/n65 ) );
  AND2_X1 \shifter_0/shift_3b_1/shift_1b_0/U3  ( .A1(
        \shifter_0/shift_3b_1/shift_1b_0/n65 ), .A2(
        \shifter_0/shift_3b_1/data1 [0]), .ZN(\shifter_0/data_3 [0]) );
  CLKBUF_X1 \shifter_0/shift_3b_1/shift_1b_0/U2  ( .A(
        \shifter_0/shift_3b_1/shift_1b_0/n64 ), .Z(
        \shifter_0/shift_3b_1/shift_1b_0/n68 ) );
  OAI21_X1 \shifter_0/shift_7b_0/U78  ( .B1(1'b0), .B2(
        \shifter_0/shift_7b_0/n79 ), .A(\shifter_0/n21 ), .ZN(
        \shifter_0/shift_7b_0/n58 ) );
  OAI21_X1 \shifter_0/shift_7b_0/U77  ( .B1(1'b0), .B2(
        \shifter_0/shift_7b_0/n80 ), .A(\shifter_0/shift_7b_0/n39 ), .ZN(
        \shifter_0/shift_7b_0/n57 ) );
  OAI21_X1 \shifter_0/shift_7b_0/U76  ( .B1(1'b0), .B2(
        \shifter_0/shift_7b_0/n78 ), .A(\shifter_0/shift_7b_0/n39 ), .ZN(
        \shifter_0/shift_7b_0/n59 ) );
  OAI22_X1 \shifter_0/shift_7b_0/U75  ( .A1(\shifter_0/shift_7b_0/n41 ), .A2(
        \shifter_0/shift_7b_0/n43 ), .B1(\shifter_0/shift_7b_0/n39 ), .B2(
        \shifter_0/shift_7b_0/n73 ), .ZN(\shifter_0/shift_7b_0/n11 ) );
  OAI22_X1 \shifter_0/shift_7b_0/U74  ( .A1(\shifter_0/shift_7b_0/n41 ), .A2(
        \shifter_0/shift_7b_0/n44 ), .B1(\shifter_0/shift_7b_0/n39 ), .B2(
        \shifter_0/shift_7b_0/n74 ), .ZN(\shifter_0/shift_7b_0/n13 ) );
  OAI22_X1 \shifter_0/shift_7b_0/U73  ( .A1(\shifter_0/shift_7b_0/n41 ), .A2(
        \shifter_0/shift_7b_0/n45 ), .B1(\shifter_0/shift_7b_0/n39 ), .B2(
        \shifter_0/shift_7b_0/n75 ), .ZN(\shifter_0/shift_7b_0/n15 ) );
  OAI22_X1 \shifter_0/shift_7b_0/U72  ( .A1(\shifter_0/shift_7b_0/n41 ), .A2(
        \shifter_0/shift_7b_0/n46 ), .B1(\shifter_0/shift_7b_0/n39 ), .B2(
        \shifter_0/shift_7b_0/n76 ), .ZN(\shifter_0/shift_7b_0/n17 ) );
  OAI22_X1 \shifter_0/shift_7b_0/U71  ( .A1(\shifter_0/shift_7b_0/n39 ), .A2(
        \shifter_0/shift_7b_0/n43 ), .B1(\shifter_0/shift_7b_0/n41 ), .B2(
        \shifter_0/shift_7b_0/n47 ), .ZN(\shifter_0/shift_7b_0/n12 ) );
  NOR2_X1 \shifter_0/shift_7b_0/U70  ( .A1(\shifter_0/shift_7b_0/n39 ), .A2(
        \shifter_0/shift_7b_0/n77 ), .ZN(\shifter_0/shift_7b_0/data1 [0]) );
  NOR2_X1 \shifter_0/shift_7b_0/U69  ( .A1(\shifter_0/shift_7b_0/n39 ), .A2(
        \shifter_0/shift_7b_0/n50 ), .ZN(\shifter_0/shift_7b_0/data1 [2]) );
  NOR2_X1 \shifter_0/shift_7b_0/U68  ( .A1(\shifter_0/shift_7b_0/n39 ), .A2(
        \shifter_0/shift_7b_0/n55 ), .ZN(\shifter_0/shift_7b_0/data1 [1]) );
  NOR2_X1 \shifter_0/shift_7b_0/U67  ( .A1(\shifter_0/shift_7b_0/n39 ), .A2(
        \shifter_0/shift_7b_0/n49 ), .ZN(\shifter_0/shift_7b_0/data1 [3]) );
  INV_X1 \shifter_0/shift_7b_0/U66  ( .A(shifted_o[3]), .ZN(
        \shifter_0/shift_7b_0/n78 ) );
  INV_X1 \shifter_0/shift_7b_0/U65  ( .A(\shifter_0/n21 ), .ZN(
        \shifter_0/shift_7b_0/n42 ) );
  INV_X1 \shifter_0/shift_7b_0/U64  ( .A(\shifter_0/n31 ), .ZN(
        \shifter_0/shift_7b_0/n80 ) );
  OAI21_X1 \shifter_0/shift_7b_0/U63  ( .B1(\shifter_0/shift_7b_0/n40 ), .B2(
        \shifter_0/shift_7b_0/n80 ), .A(\shifter_0/shift_7b_0/n57 ), .ZN(
        \shifter_0/shift_7b_0/shift1 [2]) );
  INV_X1 \shifter_0/shift_7b_0/U62  ( .A(\shifter_0/n1 ), .ZN(
        \shifter_0/shift_7b_0/n79 ) );
  OAI21_X1 \shifter_0/shift_7b_0/U61  ( .B1(\shifter_0/shift_7b_0/n40 ), .B2(
        \shifter_0/shift_7b_0/n79 ), .A(\shifter_0/shift_7b_0/n58 ), .ZN(
        \shifter_0/shift_7b_0/shift1 [1]) );
  OAI21_X1 \shifter_0/shift_7b_0/U60  ( .B1(\shifter_0/shift_7b_0/n40 ), .B2(
        \shifter_0/shift_7b_0/n78 ), .A(\shifter_0/shift_7b_0/n59 ), .ZN(
        \shifter_0/shift_7b_0/shift1 [0]) );
  INV_X1 \shifter_0/shift_7b_0/U59  ( .A(\shifter_0/data_3 [9]), .ZN(
        \shifter_0/shift_7b_0/n43 ) );
  AOI22_X1 \shifter_0/shift_7b_0/U58  ( .A1(\shifter_0/shift_7b_0/n41 ), .A2(
        \shifter_0/data_3 [31]), .B1(\shifter_0/shift_7b_0/n39 ), .B2(
        \shifter_0/data_3 [27]), .ZN(\shifter_0/shift_7b_0/n67 ) );
  INV_X1 \shifter_0/shift_7b_0/U57  ( .A(\shifter_0/shift_7b_0/n67 ), .ZN(
        \shifter_0/shift_7b_0/n21 ) );
  OAI22_X1 \shifter_0/shift_7b_0/U56  ( .A1(\shifter_0/shift_7b_0/n39 ), .A2(
        \shifter_0/shift_7b_0/n70 ), .B1(\shifter_0/shift_7b_0/n41 ), .B2(
        \shifter_0/shift_7b_0/n74 ), .ZN(\shifter_0/shift_7b_0/n36 ) );
  OAI22_X1 \shifter_0/shift_7b_0/U55  ( .A1(\shifter_0/shift_7b_0/n39 ), .A2(
        \shifter_0/shift_7b_0/n72 ), .B1(\shifter_0/shift_7b_0/n41 ), .B2(
        \shifter_0/shift_7b_0/n76 ), .ZN(\shifter_0/shift_7b_0/n38 ) );
  INV_X1 \shifter_0/shift_7b_0/U54  ( .A(\shifter_0/data_3 [11]), .ZN(
        \shifter_0/shift_7b_0/n75 ) );
  INV_X1 \shifter_0/shift_7b_0/U53  ( .A(\shifter_0/data_3 [12]), .ZN(
        \shifter_0/shift_7b_0/n74 ) );
  INV_X1 \shifter_0/shift_7b_0/U52  ( .A(\shifter_0/data_3 [13]), .ZN(
        \shifter_0/shift_7b_0/n73 ) );
  INV_X1 \shifter_0/shift_7b_0/U51  ( .A(\shifter_0/data_3 [10]), .ZN(
        \shifter_0/shift_7b_0/n76 ) );
  INV_X1 \shifter_0/shift_7b_0/U50  ( .A(\shifter_0/data_3 [8]), .ZN(
        \shifter_0/shift_7b_0/n44 ) );
  INV_X1 \shifter_0/shift_7b_0/U49  ( .A(\shifter_0/data_3 [1]), .ZN(
        \shifter_0/shift_7b_0/n55 ) );
  INV_X1 \shifter_0/shift_7b_0/U48  ( .A(\shifter_0/data_3 [7]), .ZN(
        \shifter_0/shift_7b_0/n45 ) );
  INV_X1 \shifter_0/shift_7b_0/U47  ( .A(\shifter_0/data_3 [6]), .ZN(
        \shifter_0/shift_7b_0/n46 ) );
  INV_X1 \shifter_0/shift_7b_0/U46  ( .A(\shifter_0/data_3 [2]), .ZN(
        \shifter_0/shift_7b_0/n50 ) );
  INV_X1 \shifter_0/shift_7b_0/U45  ( .A(\shifter_0/data_3 [3]), .ZN(
        \shifter_0/shift_7b_0/n49 ) );
  INV_X1 \shifter_0/shift_7b_0/U44  ( .A(\shifter_0/data_3 [5]), .ZN(
        \shifter_0/shift_7b_0/n47 ) );
  OAI22_X1 \shifter_0/shift_7b_0/U43  ( .A1(\shifter_0/shift_7b_0/n39 ), .A2(
        \shifter_0/shift_7b_0/n71 ), .B1(\shifter_0/shift_7b_0/n41 ), .B2(
        \shifter_0/shift_7b_0/n75 ), .ZN(\shifter_0/shift_7b_0/n37 ) );
  OAI22_X1 \shifter_0/shift_7b_0/U42  ( .A1(\shifter_0/shift_7b_0/n39 ), .A2(
        \shifter_0/shift_7b_0/n44 ), .B1(\shifter_0/shift_7b_0/n41 ), .B2(
        \shifter_0/shift_7b_0/n48 ), .ZN(\shifter_0/shift_7b_0/n14 ) );
  OAI22_X1 \shifter_0/shift_7b_0/U41  ( .A1(\shifter_0/shift_7b_0/n39 ), .A2(
        \shifter_0/shift_7b_0/n45 ), .B1(\shifter_0/shift_7b_0/n42 ), .B2(
        \shifter_0/shift_7b_0/n49 ), .ZN(\shifter_0/shift_7b_0/n16 ) );
  OAI22_X1 \shifter_0/shift_7b_0/U40  ( .A1(\shifter_0/shift_7b_0/n40 ), .A2(
        \shifter_0/shift_7b_0/n68 ), .B1(\shifter_0/shift_7b_0/n42 ), .B2(
        \shifter_0/shift_7b_0/n72 ), .ZN(\shifter_0/shift_7b_0/n34 ) );
  AOI22_X1 \shifter_0/shift_7b_0/U39  ( .A1(\shifter_0/shift_7b_0/n41 ), .A2(
        \shifter_0/data_3 [24]), .B1(\shifter_0/shift_7b_0/n40 ), .B2(
        \shifter_0/data_3 [20]), .ZN(\shifter_0/shift_7b_0/n60 ) );
  INV_X1 \shifter_0/shift_7b_0/U38  ( .A(\shifter_0/shift_7b_0/n60 ), .ZN(
        \shifter_0/shift_7b_0/n4 ) );
  AOI22_X1 \shifter_0/shift_7b_0/U37  ( .A1(\shifter_0/shift_7b_0/n41 ), .A2(
        \shifter_0/data_3 [25]), .B1(\shifter_0/shift_7b_0/n40 ), .B2(
        \shifter_0/data_3 [21]), .ZN(\shifter_0/shift_7b_0/n61 ) );
  INV_X1 \shifter_0/shift_7b_0/U36  ( .A(\shifter_0/shift_7b_0/n61 ), .ZN(
        \shifter_0/shift_7b_0/n5 ) );
  INV_X1 \shifter_0/shift_7b_0/U35  ( .A(\shifter_0/data_3 [4]), .ZN(
        \shifter_0/shift_7b_0/n48 ) );
  INV_X1 \shifter_0/shift_7b_0/U34  ( .A(\shifter_0/data_3 [14]), .ZN(
        \shifter_0/shift_7b_0/n72 ) );
  INV_X1 \shifter_0/shift_7b_0/U33  ( .A(\shifter_0/data_3 [17]), .ZN(
        \shifter_0/shift_7b_0/n69 ) );
  INV_X1 \shifter_0/shift_7b_0/U32  ( .A(\shifter_0/data_3 [16]), .ZN(
        \shifter_0/shift_7b_0/n70 ) );
  INV_X1 \shifter_0/shift_7b_0/U31  ( .A(\shifter_0/data_3 [15]), .ZN(
        \shifter_0/shift_7b_0/n71 ) );
  INV_X1 \shifter_0/shift_7b_0/U30  ( .A(\shifter_0/data_3 [18]), .ZN(
        \shifter_0/shift_7b_0/n68 ) );
  INV_X1 \shifter_0/shift_7b_0/U29  ( .A(\shifter_0/data_3 [19]), .ZN(
        \shifter_0/shift_7b_0/n56 ) );
  INV_X1 \shifter_0/shift_7b_0/U28  ( .A(\shifter_0/data_3 [21]), .ZN(
        \shifter_0/shift_7b_0/n53 ) );
  OAI22_X1 \shifter_0/shift_7b_0/U27  ( .A1(\shifter_0/shift_7b_0/n39 ), .A2(
        \shifter_0/shift_7b_0/n53 ), .B1(\shifter_0/shift_7b_0/n41 ), .B2(
        \shifter_0/shift_7b_0/n69 ), .ZN(\shifter_0/shift_7b_0/n31 ) );
  INV_X1 \shifter_0/shift_7b_0/U26  ( .A(\shifter_0/data_3 [20]), .ZN(
        \shifter_0/shift_7b_0/n54 ) );
  OAI22_X1 \shifter_0/shift_7b_0/U25  ( .A1(\shifter_0/shift_7b_0/n39 ), .A2(
        \shifter_0/shift_7b_0/n54 ), .B1(\shifter_0/shift_7b_0/n41 ), .B2(
        \shifter_0/shift_7b_0/n70 ), .ZN(\shifter_0/shift_7b_0/n32 ) );
  INV_X1 \shifter_0/shift_7b_0/U24  ( .A(\shifter_0/data_3 [22]), .ZN(
        \shifter_0/shift_7b_0/n52 ) );
  OAI22_X1 \shifter_0/shift_7b_0/U23  ( .A1(\shifter_0/shift_7b_0/n39 ), .A2(
        \shifter_0/shift_7b_0/n52 ), .B1(\shifter_0/shift_7b_0/n41 ), .B2(
        \shifter_0/shift_7b_0/n68 ), .ZN(\shifter_0/shift_7b_0/n30 ) );
  INV_X1 \shifter_0/shift_7b_0/U22  ( .A(\shifter_0/data_3 [23]), .ZN(
        \shifter_0/shift_7b_0/n51 ) );
  OAI22_X1 \shifter_0/shift_7b_0/U21  ( .A1(\shifter_0/shift_7b_0/n39 ), .A2(
        \shifter_0/shift_7b_0/n51 ), .B1(\shifter_0/shift_7b_0/n41 ), .B2(
        \shifter_0/shift_7b_0/n56 ), .ZN(\shifter_0/shift_7b_0/n29 ) );
  OAI22_X1 \shifter_0/shift_7b_0/U20  ( .A1(\shifter_0/shift_7b_0/n39 ), .A2(
        \shifter_0/shift_7b_0/n46 ), .B1(\shifter_0/shift_7b_0/n41 ), .B2(
        \shifter_0/shift_7b_0/n50 ), .ZN(\shifter_0/shift_7b_0/n18 ) );
  OAI22_X1 \shifter_0/shift_7b_0/U19  ( .A1(\shifter_0/shift_7b_0/n39 ), .A2(
        \shifter_0/shift_7b_0/n47 ), .B1(\shifter_0/shift_7b_0/n41 ), .B2(
        \shifter_0/shift_7b_0/n55 ), .ZN(\shifter_0/shift_7b_0/n19 ) );
  OAI22_X1 \shifter_0/shift_7b_0/U18  ( .A1(\shifter_0/shift_7b_0/n39 ), .A2(
        \shifter_0/shift_7b_0/n48 ), .B1(\shifter_0/shift_7b_0/n41 ), .B2(
        \shifter_0/shift_7b_0/n77 ), .ZN(\shifter_0/shift_7b_0/n20 ) );
  OAI22_X1 \shifter_0/shift_7b_0/U17  ( .A1(\shifter_0/shift_7b_0/n40 ), .A2(
        \shifter_0/shift_7b_0/n56 ), .B1(\shifter_0/shift_7b_0/n41 ), .B2(
        \shifter_0/shift_7b_0/n71 ), .ZN(\shifter_0/shift_7b_0/n33 ) );
  OAI22_X1 \shifter_0/shift_7b_0/U16  ( .A1(\shifter_0/shift_7b_0/n40 ), .A2(
        \shifter_0/shift_7b_0/n69 ), .B1(\shifter_0/shift_7b_0/n42 ), .B2(
        \shifter_0/shift_7b_0/n73 ), .ZN(\shifter_0/shift_7b_0/n35 ) );
  AOI22_X1 \shifter_0/shift_7b_0/U15  ( .A1(\shifter_0/shift_7b_0/n41 ), .A2(
        \shifter_0/data_3 [30]), .B1(\shifter_0/shift_7b_0/n40 ), .B2(
        \shifter_0/data_3 [26]), .ZN(\shifter_0/shift_7b_0/n66 ) );
  INV_X1 \shifter_0/shift_7b_0/U14  ( .A(\shifter_0/shift_7b_0/n66 ), .ZN(
        \shifter_0/shift_7b_0/n10 ) );
  AOI22_X1 \shifter_0/shift_7b_0/U13  ( .A1(\shifter_0/shift_7b_0/n41 ), .A2(
        \shifter_0/data_3 [26]), .B1(\shifter_0/shift_7b_0/n40 ), .B2(
        \shifter_0/data_3 [22]), .ZN(\shifter_0/shift_7b_0/n62 ) );
  INV_X1 \shifter_0/shift_7b_0/U12  ( .A(\shifter_0/shift_7b_0/n62 ), .ZN(
        \shifter_0/shift_7b_0/n6 ) );
  AOI22_X1 \shifter_0/shift_7b_0/U11  ( .A1(\shifter_0/shift_7b_0/n41 ), .A2(
        \shifter_0/data_3 [27]), .B1(\shifter_0/shift_7b_0/n40 ), .B2(
        \shifter_0/data_3 [23]), .ZN(\shifter_0/shift_7b_0/n63 ) );
  INV_X1 \shifter_0/shift_7b_0/U10  ( .A(\shifter_0/shift_7b_0/n63 ), .ZN(
        \shifter_0/shift_7b_0/n7 ) );
  AOI22_X1 \shifter_0/shift_7b_0/U9  ( .A1(\shifter_0/shift_7b_0/n41 ), .A2(
        \shifter_0/data_3 [28]), .B1(\shifter_0/shift_7b_0/n40 ), .B2(
        \shifter_0/data_3 [24]), .ZN(\shifter_0/shift_7b_0/n64 ) );
  INV_X1 \shifter_0/shift_7b_0/U8  ( .A(\shifter_0/shift_7b_0/n64 ), .ZN(
        \shifter_0/shift_7b_0/n8 ) );
  AOI22_X1 \shifter_0/shift_7b_0/U7  ( .A1(\shifter_0/shift_7b_0/n41 ), .A2(
        \shifter_0/data_3 [29]), .B1(\shifter_0/shift_7b_0/n40 ), .B2(
        \shifter_0/data_3 [25]), .ZN(\shifter_0/shift_7b_0/n65 ) );
  INV_X1 \shifter_0/shift_7b_0/U6  ( .A(\shifter_0/shift_7b_0/n65 ), .ZN(
        \shifter_0/shift_7b_0/n9 ) );
  INV_X1 \shifter_0/shift_7b_0/U5  ( .A(\shifter_0/shift_7b_0/n42 ), .ZN(
        \shifter_0/shift_7b_0/n39 ) );
  INV_X1 \shifter_0/shift_7b_0/U4  ( .A(\shifter_0/shift_7b_0/n42 ), .ZN(
        \shifter_0/shift_7b_0/n40 ) );
  INV_X1 \shifter_0/shift_7b_0/U3  ( .A(\shifter_0/data_3 [0]), .ZN(
        \shifter_0/shift_7b_0/n77 ) );
  BUF_X1 \shifter_0/shift_7b_0/U2  ( .A(\shifter_0/shift_7b_0/n42 ), .Z(
        \shifter_0/shift_7b_0/n41 ) );
  OAI21_X1 \shifter_0/shift_7b_0/shift_3b_0/U72  ( .B1(
        \shifter_0/shift_7b_0/shift1 [0]), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n39 ), .A(
        \shifter_0/shift_7b_0/shift_3b_0/n35 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/n61 ) );
  OAI22_X1 \shifter_0/shift_7b_0/shift_3b_0/U71  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/n35 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n41 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/n37 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n45 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/n5 ) );
  OAI22_X1 \shifter_0/shift_7b_0/shift_3b_0/U70  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/n35 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n70 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/n37 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n41 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/n6 ) );
  OAI22_X1 \shifter_0/shift_7b_0/shift_3b_0/U69  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/n35 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n43 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/n37 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n47 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/n9 ) );
  OAI22_X1 \shifter_0/shift_7b_0/shift_3b_0/U68  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/n35 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n71 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/n37 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n43 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/n10 ) );
  OAI22_X1 \shifter_0/shift_7b_0/shift_3b_0/U67  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/n35 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n67 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/n37 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n69 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/n32 ) );
  OAI22_X1 \shifter_0/shift_7b_0/shift_3b_0/U66  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/n35 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n69 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/n37 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n71 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/n34 ) );
  OAI22_X1 \shifter_0/shift_7b_0/shift_3b_0/U65  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/n37 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n40 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/n35 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n45 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/n7 ) );
  OAI22_X1 \shifter_0/shift_7b_0/shift_3b_0/U64  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/n37 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n42 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/n35 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n47 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/n11 ) );
  OAI22_X1 \shifter_0/shift_7b_0/shift_3b_0/U63  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/n35 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n40 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/n37 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n44 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/n8 ) );
  NOR2_X1 \shifter_0/shift_7b_0/shift_3b_0/U62  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/n35 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n60 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/data1 [1]) );
  NOR2_X1 \shifter_0/shift_7b_0/shift_3b_0/U61  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/n35 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n72 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/data1 [0]) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/U60  ( .A(
        \shifter_0/shift_7b_0/shift1 [1]), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/n38 ) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/U59  ( .A(
        \shifter_0/shift_7b_0/shift1 [2]), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/n39 ) );
  OAI21_X1 \shifter_0/shift_7b_0/shift_3b_0/U58  ( .B1(
        \shifter_0/shift_7b_0/shift_3b_0/n36 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n39 ), .A(
        \shifter_0/shift_7b_0/shift_3b_0/n61 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/shift1 ) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/U57  ( .A(\shifter_0/shift_7b_0/n36 ), .ZN(\shifter_0/shift_7b_0/shift_3b_0/n69 ) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/U56  ( .A(\shifter_0/shift_7b_0/n38 ), .ZN(\shifter_0/shift_7b_0/shift_3b_0/n71 ) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/U55  ( .A(\shifter_0/shift_7b_0/n12 ), .ZN(\shifter_0/shift_7b_0/shift_3b_0/n40 ) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/U54  ( .A(\shifter_0/shift_7b_0/n13 ), .ZN(\shifter_0/shift_7b_0/shift_3b_0/n43 ) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/U53  ( .A(\shifter_0/shift_7b_0/n11 ), .ZN(\shifter_0/shift_7b_0/shift_3b_0/n41 ) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/U52  ( .A(\shifter_0/shift_7b_0/n15 ), .ZN(\shifter_0/shift_7b_0/shift_3b_0/n45 ) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/U51  ( .A(\shifter_0/shift_7b_0/n17 ), .ZN(\shifter_0/shift_7b_0/shift_3b_0/n47 ) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/U50  ( .A(\shifter_0/shift_7b_0/n37 ), .ZN(\shifter_0/shift_7b_0/shift_3b_0/n70 ) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/U49  ( .A(\shifter_0/shift_7b_0/n14 ), .ZN(\shifter_0/shift_7b_0/shift_3b_0/n42 ) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/U48  ( .A(\shifter_0/shift_7b_0/n16 ), .ZN(\shifter_0/shift_7b_0/shift_3b_0/n44 ) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/U47  ( .A(\shifter_0/shift_7b_0/n34 ), .ZN(\shifter_0/shift_7b_0/shift_3b_0/n67 ) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/U46  ( .A(\shifter_0/shift_7b_0/n4 ), 
        .ZN(\shifter_0/shift_7b_0/shift_3b_0/n55 ) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/U45  ( .A(\shifter_0/shift_7b_0/n5 ), 
        .ZN(\shifter_0/shift_7b_0/shift_3b_0/n54 ) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/U44  ( .A(\shifter_0/shift_7b_0/n31 ), .ZN(\shifter_0/shift_7b_0/shift_3b_0/n58 ) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/U43  ( .A(\shifter_0/shift_7b_0/n32 ), .ZN(\shifter_0/shift_7b_0/shift_3b_0/n59 ) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/U42  ( .A(\shifter_0/shift_7b_0/n30 ), .ZN(\shifter_0/shift_7b_0/shift_3b_0/n57 ) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/U41  ( .A(\shifter_0/shift_7b_0/n29 ), .ZN(\shifter_0/shift_7b_0/shift_3b_0/n56 ) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/U40  ( .A(\shifter_0/shift_7b_0/n18 ), .ZN(\shifter_0/shift_7b_0/shift_3b_0/n46 ) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/U39  ( .A(\shifter_0/shift_7b_0/n19 ), .ZN(\shifter_0/shift_7b_0/shift_3b_0/n48 ) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/U38  ( .A(\shifter_0/shift_7b_0/n20 ), .ZN(\shifter_0/shift_7b_0/shift_3b_0/n49 ) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/U37  ( .A(\shifter_0/shift_7b_0/n33 ), .ZN(\shifter_0/shift_7b_0/shift_3b_0/n66 ) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/U36  ( .A(\shifter_0/shift_7b_0/n35 ), .ZN(\shifter_0/shift_7b_0/shift_3b_0/n68 ) );
  AOI22_X1 \shifter_0/shift_7b_0/shift_3b_0/U35  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/n37 ), .A2(\shifter_0/shift_7b_0/n8 ), 
        .B1(\shifter_0/shift_7b_0/shift_3b_0/n36 ), .B2(
        \shifter_0/shift_7b_0/n6 ), .ZN(\shifter_0/shift_7b_0/shift_3b_0/n62 )
         );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/U34  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/n62 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/n2 ) );
  AOI22_X1 \shifter_0/shift_7b_0/shift_3b_0/U33  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/n37 ), .A2(\shifter_0/shift_7b_0/n10 ), .B1(\shifter_0/shift_7b_0/shift_3b_0/n36 ), .B2(\shifter_0/shift_7b_0/n8 ), 
        .ZN(\shifter_0/shift_7b_0/shift_3b_0/n64 ) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/U32  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/n64 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/n4 ) );
  AOI22_X1 \shifter_0/shift_7b_0/shift_3b_0/U31  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/n37 ), .A2(\shifter_0/shift_7b_0/n9 ), 
        .B1(\shifter_0/shift_7b_0/shift_3b_0/n36 ), .B2(
        \shifter_0/shift_7b_0/n7 ), .ZN(\shifter_0/shift_7b_0/shift_3b_0/n63 )
         );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/U30  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/n63 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/n3 ) );
  AOI22_X1 \shifter_0/shift_7b_0/shift_3b_0/U29  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/n37 ), .A2(\shifter_0/shift_7b_0/n21 ), .B1(\shifter_0/shift_7b_0/shift_3b_0/n36 ), .B2(\shifter_0/shift_7b_0/n9 ), 
        .ZN(\shifter_0/shift_7b_0/shift_3b_0/n65 ) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/U28  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/n65 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/n18 ) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/U27  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/n38 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/n35 ) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/U26  ( .A(\shifter_0/shift_7b_0/n6 ), 
        .ZN(\shifter_0/shift_7b_0/shift_3b_0/n53 ) );
  OAI22_X1 \shifter_0/shift_7b_0/shift_3b_0/U25  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/n36 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n53 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/n38 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n55 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/n24 ) );
  OAI22_X1 \shifter_0/shift_7b_0/shift_3b_0/U24  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/n36 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n59 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/n37 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n67 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/n30 ) );
  OAI22_X1 \shifter_0/shift_7b_0/shift_3b_0/U23  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/n36 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n56 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/n37 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n58 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/n27 ) );
  OAI22_X1 \shifter_0/shift_7b_0/shift_3b_0/U22  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/n36 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n57 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/n37 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n59 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/n28 ) );
  OAI22_X1 \shifter_0/shift_7b_0/shift_3b_0/U21  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/n36 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n58 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/n37 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n66 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/n29 ) );
  OAI22_X1 \shifter_0/shift_7b_0/shift_3b_0/U20  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/n36 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n55 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/n37 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n57 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/n26 ) );
  OAI22_X1 \shifter_0/shift_7b_0/shift_3b_0/U19  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/n36 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n54 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/n37 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n56 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/n25 ) );
  OAI22_X1 \shifter_0/shift_7b_0/shift_3b_0/U18  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/n36 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n68 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/n37 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n70 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/n33 ) );
  OAI22_X1 \shifter_0/shift_7b_0/shift_3b_0/U17  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/n36 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n66 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/n37 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n68 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/n31 ) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/U16  ( .A(\shifter_0/shift_7b_0/n7 ), 
        .ZN(\shifter_0/shift_7b_0/shift_3b_0/n52 ) );
  OAI22_X1 \shifter_0/shift_7b_0/shift_3b_0/U15  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/n36 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n52 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/n38 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n54 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/n23 ) );
  OAI22_X1 \shifter_0/shift_7b_0/shift_3b_0/U14  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/n36 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n42 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/n37 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n46 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/n12 ) );
  OAI22_X1 \shifter_0/shift_7b_0/shift_3b_0/U13  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/n36 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n51 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/n37 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n72 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/n20 ) );
  OAI22_X1 \shifter_0/shift_7b_0/shift_3b_0/U12  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/n36 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n50 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/n38 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n60 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/n17 ) );
  OAI22_X1 \shifter_0/shift_7b_0/shift_3b_0/U11  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/n36 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n48 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/n37 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n50 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/n15 ) );
  OAI22_X1 \shifter_0/shift_7b_0/shift_3b_0/U10  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/n36 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n44 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/n37 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n48 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/n13 ) );
  OAI22_X1 \shifter_0/shift_7b_0/shift_3b_0/U9  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/n36 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n49 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/n38 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n51 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/n16 ) );
  OAI22_X1 \shifter_0/shift_7b_0/shift_3b_0/U8  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/n36 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n46 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/n38 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n49 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/n14 ) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/U7  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/n38 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/n36 ) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/U6  ( .A(
        \shifter_0/shift_7b_0/data1 [0]), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/n72 ) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/U5  ( .A(
        \shifter_0/shift_7b_0/data1 [1]), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/n60 ) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/U4  ( .A(
        \shifter_0/shift_7b_0/data1 [3]), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/n50 ) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/U3  ( .A(
        \shifter_0/shift_7b_0/data1 [2]), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/n51 ) );
  BUF_X1 \shifter_0/shift_7b_0/shift_3b_0/U2  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/n38 ), .Z(
        \shifter_0/shift_7b_0/shift_3b_0/n37 ) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U68  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n67 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n66 ) );
  AOI22_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U67  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n67 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n8 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n66 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n11 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n63 ) );
  AOI22_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U66  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n66 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n9 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n64 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n7 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n61 ) );
  AOI22_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U65  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n66 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n5 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n64 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n9 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n60 ) );
  AOI22_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U64  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n66 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n10 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n64 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n5 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n59 ) );
  AOI22_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U63  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n66 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n6 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n64 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n10 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n58 ) );
  AOI22_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U62  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n66 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n34 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n64 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n6 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n57 ) );
  AOI22_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U61  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n66 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n7 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n64 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n11 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n62 ) );
  AND2_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U60  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n66 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/data1 [0]), .ZN(sdata_o[0]) );
  AOI22_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U59  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n65 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/data1 [1]), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n64 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/data1 [0]), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n53 ) );
  AOI22_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U58  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n66 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n32 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n64 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n33 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n55 ) );
  AOI22_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U57  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n65 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n33 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n64 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n34 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n56 ) );
  AOI22_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U56  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n65 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n31 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n64 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n32 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n54 ) );
  AOI22_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U55  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n66 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n30 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n64 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n31 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n52 ) );
  AOI22_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U54  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n65 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n29 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n64 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n30 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n51 ) );
  AOI22_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U53  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n66 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n28 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n64 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n29 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n50 ) );
  AOI22_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U52  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n65 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n27 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n64 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n28 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n49 ) );
  AOI22_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U51  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n66 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n26 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n64 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n27 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n48 ) );
  AOI22_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U50  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n66 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n25 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n64 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n26 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n47 ) );
  AOI22_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U49  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n65 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n24 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n64 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n25 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n46 ) );
  AOI22_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U48  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n66 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n23 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n64 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n24 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n45 ) );
  AOI22_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U47  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n65 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n18 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n64 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n4 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n40 ) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U46  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n40 ), .ZN(sdata_o[31]) );
  BUF_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U45  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/shift1 ), .Z(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n67 ) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U44  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n45 ), .ZN(sdata_o[27]) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U43  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n51 ), .ZN(sdata_o[21]) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U42  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n48 ), .ZN(sdata_o[24]) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U41  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n49 ), .ZN(sdata_o[23]) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U40  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n50 ), .ZN(sdata_o[22]) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U39  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n47 ), .ZN(sdata_o[25]) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U38  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n46 ), .ZN(sdata_o[26]) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U37  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n55 ), .ZN(sdata_o[18]) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U36  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n52 ), .ZN(sdata_o[20]) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U35  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n53 ), .ZN(sdata_o[1]) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U34  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n56 ), .ZN(sdata_o[17]) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U33  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n54 ), .ZN(sdata_o[19]) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U32  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n61 ), .ZN(sdata_o[12]) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U31  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n59 ), .ZN(sdata_o[14]) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U30  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n60 ), .ZN(sdata_o[13]) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U29  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n58 ), .ZN(sdata_o[15]) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U28  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n62 ), .ZN(sdata_o[11]) );
  AOI22_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U27  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n65 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n14 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n64 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n15 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n36 ) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U26  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n36 ), .ZN(sdata_o[6]) );
  AOI22_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U25  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n65 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n12 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n67 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n13 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n34 ) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U24  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n34 ), .ZN(sdata_o[8]) );
  AOI22_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U23  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n65 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n13 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n67 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n14 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n35 ) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U22  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n35 ), .ZN(sdata_o[7]) );
  AOI22_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U21  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n65 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n3 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n64 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n2 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n43 ) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U20  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n43 ), .ZN(sdata_o[29]) );
  AOI22_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U19  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n65 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n4 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n64 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n3 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n41 ) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U18  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n41 ), .ZN(sdata_o[30]) );
  AOI22_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U17  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n65 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n17 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n64 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n20 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n39 ) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U16  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n39 ), .ZN(sdata_o[3]) );
  AOI22_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U15  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n65 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n20 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/shift1 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/data1 [1]), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n42 ) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U14  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n42 ), .ZN(sdata_o[2]) );
  AOI22_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U13  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n65 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n16 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n64 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n17 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n38 ) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U12  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n38 ), .ZN(sdata_o[4]) );
  AOI22_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U11  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n65 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n15 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n64 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n16 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n37 ) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U10  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n37 ), .ZN(sdata_o[5]) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U9  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n63 ), .ZN(sdata_o[10]) );
  AOI22_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U8  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n65 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n2 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/shift1 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/n23 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n44 ) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U7  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n44 ), .ZN(sdata_o[28]) );
  AOI22_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U6  ( .A1(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n65 ), .A2(
        \shifter_0/shift_7b_0/shift_3b_0/n8 ), .B1(
        \shifter_0/shift_7b_0/shift_3b_0/n12 ), .B2(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n67 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n33 ) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U5  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n33 ), .ZN(sdata_o[9]) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U4  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n57 ), .ZN(sdata_o[16]) );
  INV_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U3  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n67 ), .ZN(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n65 ) );
  BUF_X1 \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/U2  ( .A(
        \shifter_0/shift_7b_0/shift_3b_0/shift1 ), .Z(
        \shifter_0/shift_7b_0/shift_3b_0/shift_1b_0/n64 ) );
  XOR2_X1 \adder_0/U32  ( .A(reg_carry), .B(\adder_0/P0[0] ), .Z(sum[0]) );
  XOR2_X1 \adder_0/U31  ( .A(\adder_0/P0[10] ), .B(\adder_0/G6_9 ), .Z(sum[10]) );
  XOR2_X1 \adder_0/U30  ( .A(\adder_0/P0[11] ), .B(\adder_0/G4[5] ), .Z(
        sum[11]) );
  XOR2_X1 \adder_0/U29  ( .A(\adder_0/P0[12] ), .B(\adder_0/G6_11 ), .Z(
        sum[12]) );
  XOR2_X1 \adder_0/U28  ( .A(\adder_0/P0[13] ), .B(\adder_0/G4[6] ), .Z(
        sum[13]) );
  XOR2_X1 \adder_0/U27  ( .A(\adder_0/P0[14] ), .B(\adder_0/G6_13 ), .Z(
        sum[14]) );
  XOR2_X1 \adder_0/U26  ( .A(\adder_0/P0[15] ), .B(\adder_0/G4[7] ), .Z(
        sum[15]) );
  XOR2_X1 \adder_0/U25  ( .A(\adder_0/P0[16] ), .B(\adder_0/G6_15 ), .Z(
        sum[16]) );
  XOR2_X1 \adder_0/U24  ( .A(\adder_0/P0[17] ), .B(\adder_0/G5[8] ), .Z(
        sum[17]) );
  XOR2_X1 \adder_0/U23  ( .A(\adder_0/P0[18] ), .B(\adder_0/G6_17 ), .Z(
        sum[18]) );
  XOR2_X1 \adder_0/U22  ( .A(\adder_0/P0[19] ), .B(\adder_0/G5[9] ), .Z(
        sum[19]) );
  XOR2_X1 \adder_0/U21  ( .A(\adder_0/P0[1] ), .B(\adder_0/G1[0] ), .Z(sum[1])
         );
  XOR2_X1 \adder_0/U20  ( .A(\adder_0/P0[20] ), .B(\adder_0/G6_19 ), .Z(
        sum[20]) );
  XOR2_X1 \adder_0/U19  ( .A(\adder_0/P0[21] ), .B(\adder_0/G5[10] ), .Z(
        sum[21]) );
  XOR2_X1 \adder_0/U18  ( .A(\adder_0/P0[22] ), .B(\adder_0/G6_21 ), .Z(
        sum[22]) );
  XOR2_X1 \adder_0/U17  ( .A(\adder_0/P0[23] ), .B(\adder_0/G5[11] ), .Z(
        sum[23]) );
  XOR2_X1 \adder_0/U16  ( .A(\adder_0/P0[24] ), .B(\adder_0/G6_23 ), .Z(
        sum[24]) );
  XOR2_X1 \adder_0/U15  ( .A(\adder_0/P0[25] ), .B(\adder_0/G5[12] ), .Z(
        sum[25]) );
  XOR2_X1 \adder_0/U14  ( .A(\adder_0/P0[26] ), .B(\adder_0/G6_25 ), .Z(
        sum[26]) );
  XOR2_X1 \adder_0/U13  ( .A(\adder_0/P0[27] ), .B(\adder_0/G5[13] ), .Z(
        sum[27]) );
  XOR2_X1 \adder_0/U12  ( .A(\adder_0/P0[28] ), .B(\adder_0/G6_27 ), .Z(
        sum[28]) );
  XOR2_X1 \adder_0/U11  ( .A(\adder_0/P0[29] ), .B(\adder_0/G5[14] ), .Z(
        sum[29]) );
  XOR2_X1 \adder_0/U10  ( .A(\adder_0/P0[2] ), .B(\adder_0/G6_1 ), .Z(sum[2])
         );
  XOR2_X1 \adder_0/U9  ( .A(\adder_0/P0[30] ), .B(\adder_0/G6_29_ ), .Z(
        sum[30]) );
  XOR2_X1 \adder_0/U8  ( .A(\adder_0/P0[31] ), .B(\adder_0/G5[15] ), .Z(
        sum[31]) );
  XOR2_X1 \adder_0/U7  ( .A(\adder_0/P0[3] ), .B(\adder_0/G2[1] ), .Z(sum[3])
         );
  XOR2_X1 \adder_0/U6  ( .A(\adder_0/P0[4] ), .B(\adder_0/G6_3 ), .Z(sum[4])
         );
  XOR2_X1 \adder_0/U5  ( .A(\adder_0/P0[5] ), .B(\adder_0/G3[2] ), .Z(sum[5])
         );
  XOR2_X1 \adder_0/U4  ( .A(\adder_0/P0[6] ), .B(\adder_0/G6_5 ), .Z(sum[6])
         );
  XOR2_X1 \adder_0/U3  ( .A(\adder_0/P0[7] ), .B(\adder_0/G3[3] ), .Z(sum[7])
         );
  XOR2_X1 \adder_0/U2  ( .A(\adder_0/P0[8] ), .B(\adder_0/G6_7 ), .Z(sum[8])
         );
  XOR2_X1 \adder_0/U1  ( .A(\adder_0/P0[9] ), .B(\adder_0/G4[4] ), .Z(sum[9])
         );
  AND2_X1 \adder_0/operator_A_0/U1  ( .A1(reg_b[0]), .A2(reg_a[0]), .ZN(
        \adder_0/G0[0] ) );
  XOR2_X1 \adder_0/operator_A_0/U2  ( .A(reg_b[0]), .B(reg_a[0]), .Z(
        \adder_0/P0[0] ) );
  AND2_X1 \adder_0/operator_A_1/U1  ( .A1(reg_b[1]), .A2(reg_a[1]), .ZN(
        \adder_0/G0[1] ) );
  XOR2_X1 \adder_0/operator_A_1/U2  ( .A(reg_b[1]), .B(reg_a[1]), .Z(
        \adder_0/P0[1] ) );
  AND2_X1 \adder_0/operator_A_2/U1  ( .A1(reg_b[2]), .A2(reg_a[2]), .ZN(
        \adder_0/G0[2] ) );
  XOR2_X1 \adder_0/operator_A_2/U2  ( .A(reg_b[2]), .B(reg_a[2]), .Z(
        \adder_0/P0[2] ) );
  AND2_X1 \adder_0/operator_A_3/U1  ( .A1(reg_b[3]), .A2(reg_a[3]), .ZN(
        \adder_0/G0[3] ) );
  XOR2_X1 \adder_0/operator_A_3/U2  ( .A(reg_b[3]), .B(reg_a[3]), .Z(
        \adder_0/P0[3] ) );
  AND2_X1 \adder_0/operator_A_4/U1  ( .A1(reg_b[4]), .A2(reg_a[4]), .ZN(
        \adder_0/G0[4] ) );
  XOR2_X1 \adder_0/operator_A_4/U2  ( .A(reg_b[4]), .B(reg_a[4]), .Z(
        \adder_0/P0[4] ) );
  AND2_X1 \adder_0/operator_A_5/U1  ( .A1(reg_b[5]), .A2(reg_a[5]), .ZN(
        \adder_0/G0[5] ) );
  XOR2_X1 \adder_0/operator_A_5/U2  ( .A(reg_b[5]), .B(reg_a[5]), .Z(
        \adder_0/P0[5] ) );
  AND2_X1 \adder_0/operator_A_6/U1  ( .A1(reg_b[6]), .A2(reg_a[6]), .ZN(
        \adder_0/G0[6] ) );
  XOR2_X1 \adder_0/operator_A_6/U2  ( .A(reg_b[6]), .B(reg_a[6]), .Z(
        \adder_0/P0[6] ) );
  AND2_X1 \adder_0/operator_A_7/U1  ( .A1(reg_b[7]), .A2(reg_a[7]), .ZN(
        \adder_0/G0[7] ) );
  XOR2_X1 \adder_0/operator_A_7/U2  ( .A(reg_b[7]), .B(reg_a[7]), .Z(
        \adder_0/P0[7] ) );
  AND2_X1 \adder_0/operator_A_8/U1  ( .A1(reg_b[8]), .A2(reg_a[8]), .ZN(
        \adder_0/G0[8] ) );
  XOR2_X1 \adder_0/operator_A_8/U2  ( .A(reg_b[8]), .B(reg_a[8]), .Z(
        \adder_0/P0[8] ) );
  AND2_X1 \adder_0/operator_A_9/U1  ( .A1(reg_b[9]), .A2(reg_a[9]), .ZN(
        \adder_0/G0[9] ) );
  XOR2_X1 \adder_0/operator_A_9/U2  ( .A(reg_b[9]), .B(reg_a[9]), .Z(
        \adder_0/P0[9] ) );
  AND2_X1 \adder_0/operator_A_10/U1  ( .A1(reg_b[10]), .A2(reg_a[10]), .ZN(
        \adder_0/G0[10] ) );
  XOR2_X1 \adder_0/operator_A_10/U2  ( .A(reg_b[10]), .B(reg_a[10]), .Z(
        \adder_0/P0[10] ) );
  AND2_X1 \adder_0/operator_A_11/U1  ( .A1(reg_b[11]), .A2(reg_a[11]), .ZN(
        \adder_0/G0[11] ) );
  XOR2_X1 \adder_0/operator_A_11/U2  ( .A(reg_b[11]), .B(reg_a[11]), .Z(
        \adder_0/P0[11] ) );
  AND2_X1 \adder_0/operator_A_12/U1  ( .A1(reg_b[12]), .A2(reg_a[12]), .ZN(
        \adder_0/G0[12] ) );
  XOR2_X1 \adder_0/operator_A_12/U2  ( .A(reg_b[12]), .B(reg_a[12]), .Z(
        \adder_0/P0[12] ) );
  AND2_X1 \adder_0/operator_A_13/U1  ( .A1(reg_b[13]), .A2(reg_a[13]), .ZN(
        \adder_0/G0[13] ) );
  XOR2_X1 \adder_0/operator_A_13/U2  ( .A(reg_b[13]), .B(reg_a[13]), .Z(
        \adder_0/P0[13] ) );
  AND2_X1 \adder_0/operator_A_14/U1  ( .A1(reg_b[14]), .A2(reg_a[14]), .ZN(
        \adder_0/G0[14] ) );
  XOR2_X1 \adder_0/operator_A_14/U2  ( .A(reg_b[14]), .B(reg_a[14]), .Z(
        \adder_0/P0[14] ) );
  AND2_X1 \adder_0/operator_A_15/U1  ( .A1(reg_b[15]), .A2(reg_a[15]), .ZN(
        \adder_0/G0[15] ) );
  XOR2_X1 \adder_0/operator_A_15/U2  ( .A(reg_b[15]), .B(reg_a[15]), .Z(
        \adder_0/P0[15] ) );
  AND2_X1 \adder_0/operator_A_16/U1  ( .A1(reg_b[16]), .A2(reg_a[16]), .ZN(
        \adder_0/G0[16] ) );
  XOR2_X1 \adder_0/operator_A_16/U2  ( .A(reg_b[16]), .B(reg_a[16]), .Z(
        \adder_0/P0[16] ) );
  AND2_X1 \adder_0/operator_A_17/U1  ( .A1(reg_b[17]), .A2(reg_a[17]), .ZN(
        \adder_0/G0[17] ) );
  XOR2_X1 \adder_0/operator_A_17/U2  ( .A(reg_b[17]), .B(reg_a[17]), .Z(
        \adder_0/P0[17] ) );
  AND2_X1 \adder_0/operator_A_18/U1  ( .A1(reg_b[18]), .A2(reg_a[18]), .ZN(
        \adder_0/G0[18] ) );
  XOR2_X1 \adder_0/operator_A_18/U2  ( .A(reg_b[18]), .B(reg_a[18]), .Z(
        \adder_0/P0[18] ) );
  AND2_X1 \adder_0/operator_A_19/U1  ( .A1(reg_b[19]), .A2(reg_a[19]), .ZN(
        \adder_0/G0[19] ) );
  XOR2_X1 \adder_0/operator_A_19/U2  ( .A(reg_b[19]), .B(reg_a[19]), .Z(
        \adder_0/P0[19] ) );
  AND2_X1 \adder_0/operator_A_20/U1  ( .A1(reg_b[20]), .A2(reg_a[20]), .ZN(
        \adder_0/G0[20] ) );
  XOR2_X1 \adder_0/operator_A_20/U2  ( .A(reg_b[20]), .B(reg_a[20]), .Z(
        \adder_0/P0[20] ) );
  AND2_X1 \adder_0/operator_A_21/U1  ( .A1(reg_b[21]), .A2(reg_a[21]), .ZN(
        \adder_0/G0[21] ) );
  XOR2_X1 \adder_0/operator_A_21/U2  ( .A(reg_b[21]), .B(reg_a[21]), .Z(
        \adder_0/P0[21] ) );
  AND2_X1 \adder_0/operator_A_22/U1  ( .A1(reg_b[22]), .A2(reg_a[22]), .ZN(
        \adder_0/G0[22] ) );
  XOR2_X1 \adder_0/operator_A_22/U2  ( .A(reg_b[22]), .B(reg_a[22]), .Z(
        \adder_0/P0[22] ) );
  AND2_X1 \adder_0/operator_A_23/U1  ( .A1(reg_b[23]), .A2(reg_a[23]), .ZN(
        \adder_0/G0[23] ) );
  XOR2_X1 \adder_0/operator_A_23/U2  ( .A(reg_b[23]), .B(reg_a[23]), .Z(
        \adder_0/P0[23] ) );
  AND2_X1 \adder_0/operator_A_24/U1  ( .A1(reg_b[24]), .A2(reg_a[24]), .ZN(
        \adder_0/G0[24] ) );
  XOR2_X1 \adder_0/operator_A_24/U2  ( .A(reg_b[24]), .B(reg_a[24]), .Z(
        \adder_0/P0[24] ) );
  AND2_X1 \adder_0/operator_A_25/U1  ( .A1(reg_b[25]), .A2(reg_a[25]), .ZN(
        \adder_0/G0[25] ) );
  XOR2_X1 \adder_0/operator_A_25/U2  ( .A(reg_b[25]), .B(reg_a[25]), .Z(
        \adder_0/P0[25] ) );
  AND2_X1 \adder_0/operator_A_26/U1  ( .A1(reg_b[26]), .A2(reg_a[26]), .ZN(
        \adder_0/G0[26] ) );
  XOR2_X1 \adder_0/operator_A_26/U2  ( .A(reg_b[26]), .B(reg_a[26]), .Z(
        \adder_0/P0[26] ) );
  AND2_X1 \adder_0/operator_A_27/U1  ( .A1(reg_b[27]), .A2(reg_a[27]), .ZN(
        \adder_0/G0[27] ) );
  XOR2_X1 \adder_0/operator_A_27/U2  ( .A(reg_b[27]), .B(reg_a[27]), .Z(
        \adder_0/P0[27] ) );
  AND2_X1 \adder_0/operator_A_28/U1  ( .A1(reg_b[28]), .A2(reg_a[28]), .ZN(
        \adder_0/G0[28] ) );
  XOR2_X1 \adder_0/operator_A_28/U2  ( .A(reg_b[28]), .B(reg_a[28]), .Z(
        \adder_0/P0[28] ) );
  AND2_X1 \adder_0/operator_A_29/U1  ( .A1(reg_b[29]), .A2(reg_a[29]), .ZN(
        \adder_0/G0[29] ) );
  XOR2_X1 \adder_0/operator_A_29/U2  ( .A(reg_b[29]), .B(reg_a[29]), .Z(
        \adder_0/P0[29] ) );
  AND2_X1 \adder_0/operator_A_30/U1  ( .A1(reg_b[30]), .A2(reg_a[30]), .ZN(
        \adder_0/G0[30] ) );
  XOR2_X1 \adder_0/operator_A_30/U2  ( .A(reg_b[30]), .B(reg_a[30]), .Z(
        \adder_0/P0[30] ) );
  AND2_X1 \adder_0/operator_A_31/U1  ( .A1(reg_b[31]), .A2(reg_a[31]), .ZN(
        \adder_0/G0[31] ) );
  XOR2_X1 \adder_0/operator_A_31/U2  ( .A(reg_b[31]), .B(reg_a[31]), .Z(
        \adder_0/P0[31] ) );
  AOI21_X1 \adder_0/operator_C_stage_1_0/U2  ( .B1(\adder_0/P0[0] ), .B2(
        reg_carry), .A(\adder_0/G0[0] ), .ZN(\adder_0/operator_C_stage_1_0/n2 ) );
  INV_X1 \adder_0/operator_C_stage_1_0/U1  ( .A(
        \adder_0/operator_C_stage_1_0/n2 ), .ZN(\adder_0/G1[0] ) );
  AOI21_X1 \adder_0/operator_B_stage_1_1/U3  ( .B1(\adder_0/G0[1] ), .B2(
        \adder_0/P0[2] ), .A(\adder_0/G0[2] ), .ZN(
        \adder_0/operator_B_stage_1_1/n2 ) );
  INV_X1 \adder_0/operator_B_stage_1_1/U2  ( .A(
        \adder_0/operator_B_stage_1_1/n2 ), .ZN(\adder_0/G1[1] ) );
  AND2_X1 \adder_0/operator_B_stage_1_1/U1  ( .A1(\adder_0/P0[1] ), .A2(
        \adder_0/P0[2] ), .ZN(\adder_0/P1[1] ) );
  AOI21_X1 \adder_0/operator_B_stage_1_2/U3  ( .B1(\adder_0/G0[3] ), .B2(
        \adder_0/P0[4] ), .A(\adder_0/G0[4] ), .ZN(
        \adder_0/operator_B_stage_1_2/n3 ) );
  INV_X1 \adder_0/operator_B_stage_1_2/U2  ( .A(
        \adder_0/operator_B_stage_1_2/n3 ), .ZN(\adder_0/G1[2] ) );
  AND2_X1 \adder_0/operator_B_stage_1_2/U1  ( .A1(\adder_0/P0[3] ), .A2(
        \adder_0/P0[4] ), .ZN(\adder_0/P1[2] ) );
  AOI21_X1 \adder_0/operator_B_stage_1_3/U3  ( .B1(\adder_0/G0[5] ), .B2(
        \adder_0/P0[6] ), .A(\adder_0/G0[6] ), .ZN(
        \adder_0/operator_B_stage_1_3/n3 ) );
  INV_X1 \adder_0/operator_B_stage_1_3/U2  ( .A(
        \adder_0/operator_B_stage_1_3/n3 ), .ZN(\adder_0/G1[3] ) );
  AND2_X1 \adder_0/operator_B_stage_1_3/U1  ( .A1(\adder_0/P0[5] ), .A2(
        \adder_0/P0[6] ), .ZN(\adder_0/P1[3] ) );
  AOI21_X1 \adder_0/operator_B_stage_1_4/U3  ( .B1(\adder_0/G0[7] ), .B2(
        \adder_0/P0[8] ), .A(\adder_0/G0[8] ), .ZN(
        \adder_0/operator_B_stage_1_4/n3 ) );
  INV_X1 \adder_0/operator_B_stage_1_4/U2  ( .A(
        \adder_0/operator_B_stage_1_4/n3 ), .ZN(\adder_0/G1[4] ) );
  AND2_X1 \adder_0/operator_B_stage_1_4/U1  ( .A1(\adder_0/P0[7] ), .A2(
        \adder_0/P0[8] ), .ZN(\adder_0/P1[4] ) );
  AOI21_X1 \adder_0/operator_B_stage_1_5/U3  ( .B1(\adder_0/G0[9] ), .B2(
        \adder_0/P0[10] ), .A(\adder_0/G0[10] ), .ZN(
        \adder_0/operator_B_stage_1_5/n3 ) );
  INV_X1 \adder_0/operator_B_stage_1_5/U2  ( .A(
        \adder_0/operator_B_stage_1_5/n3 ), .ZN(\adder_0/G1[5] ) );
  AND2_X1 \adder_0/operator_B_stage_1_5/U1  ( .A1(\adder_0/P0[9] ), .A2(
        \adder_0/P0[10] ), .ZN(\adder_0/P1[5] ) );
  AOI21_X1 \adder_0/operator_B_stage_1_6/U3  ( .B1(\adder_0/G0[11] ), .B2(
        \adder_0/P0[12] ), .A(\adder_0/G0[12] ), .ZN(
        \adder_0/operator_B_stage_1_6/n3 ) );
  INV_X1 \adder_0/operator_B_stage_1_6/U2  ( .A(
        \adder_0/operator_B_stage_1_6/n3 ), .ZN(\adder_0/G1[6] ) );
  AND2_X1 \adder_0/operator_B_stage_1_6/U1  ( .A1(\adder_0/P0[11] ), .A2(
        \adder_0/P0[12] ), .ZN(\adder_0/P1[6] ) );
  AOI21_X1 \adder_0/operator_B_stage_1_7/U3  ( .B1(\adder_0/G0[13] ), .B2(
        \adder_0/P0[14] ), .A(\adder_0/G0[14] ), .ZN(
        \adder_0/operator_B_stage_1_7/n3 ) );
  INV_X1 \adder_0/operator_B_stage_1_7/U2  ( .A(
        \adder_0/operator_B_stage_1_7/n3 ), .ZN(\adder_0/G1[7] ) );
  AND2_X1 \adder_0/operator_B_stage_1_7/U1  ( .A1(\adder_0/P0[13] ), .A2(
        \adder_0/P0[14] ), .ZN(\adder_0/P1[7] ) );
  AOI21_X1 \adder_0/operator_B_stage_1_8/U3  ( .B1(\adder_0/G0[15] ), .B2(
        \adder_0/P0[16] ), .A(\adder_0/G0[16] ), .ZN(
        \adder_0/operator_B_stage_1_8/n3 ) );
  INV_X1 \adder_0/operator_B_stage_1_8/U2  ( .A(
        \adder_0/operator_B_stage_1_8/n3 ), .ZN(\adder_0/G1[8] ) );
  AND2_X1 \adder_0/operator_B_stage_1_8/U1  ( .A1(\adder_0/P0[15] ), .A2(
        \adder_0/P0[16] ), .ZN(\adder_0/P1[8] ) );
  AOI21_X1 \adder_0/operator_B_stage_1_9/U3  ( .B1(\adder_0/G0[17] ), .B2(
        \adder_0/P0[18] ), .A(\adder_0/G0[18] ), .ZN(
        \adder_0/operator_B_stage_1_9/n3 ) );
  INV_X1 \adder_0/operator_B_stage_1_9/U2  ( .A(
        \adder_0/operator_B_stage_1_9/n3 ), .ZN(\adder_0/G1[9] ) );
  AND2_X1 \adder_0/operator_B_stage_1_9/U1  ( .A1(\adder_0/P0[17] ), .A2(
        \adder_0/P0[18] ), .ZN(\adder_0/P1[9] ) );
  AOI21_X1 \adder_0/operator_B_stage_1_10/U3  ( .B1(\adder_0/G0[19] ), .B2(
        \adder_0/P0[20] ), .A(\adder_0/G0[20] ), .ZN(
        \adder_0/operator_B_stage_1_10/n3 ) );
  INV_X1 \adder_0/operator_B_stage_1_10/U2  ( .A(
        \adder_0/operator_B_stage_1_10/n3 ), .ZN(\adder_0/G1[10] ) );
  AND2_X1 \adder_0/operator_B_stage_1_10/U1  ( .A1(\adder_0/P0[19] ), .A2(
        \adder_0/P0[20] ), .ZN(\adder_0/P1[10] ) );
  AOI21_X1 \adder_0/operator_B_stage_1_11/U3  ( .B1(\adder_0/G0[21] ), .B2(
        \adder_0/P0[22] ), .A(\adder_0/G0[22] ), .ZN(
        \adder_0/operator_B_stage_1_11/n3 ) );
  INV_X1 \adder_0/operator_B_stage_1_11/U2  ( .A(
        \adder_0/operator_B_stage_1_11/n3 ), .ZN(\adder_0/G1[11] ) );
  AND2_X1 \adder_0/operator_B_stage_1_11/U1  ( .A1(\adder_0/P0[21] ), .A2(
        \adder_0/P0[22] ), .ZN(\adder_0/P1[11] ) );
  AOI21_X1 \adder_0/operator_B_stage_1_12/U3  ( .B1(\adder_0/G0[23] ), .B2(
        \adder_0/P0[24] ), .A(\adder_0/G0[24] ), .ZN(
        \adder_0/operator_B_stage_1_12/n3 ) );
  INV_X1 \adder_0/operator_B_stage_1_12/U2  ( .A(
        \adder_0/operator_B_stage_1_12/n3 ), .ZN(\adder_0/G1[12] ) );
  AND2_X1 \adder_0/operator_B_stage_1_12/U1  ( .A1(\adder_0/P0[23] ), .A2(
        \adder_0/P0[24] ), .ZN(\adder_0/P1[12] ) );
  AOI21_X1 \adder_0/operator_B_stage_1_13/U3  ( .B1(\adder_0/G0[25] ), .B2(
        \adder_0/P0[26] ), .A(\adder_0/G0[26] ), .ZN(
        \adder_0/operator_B_stage_1_13/n3 ) );
  INV_X1 \adder_0/operator_B_stage_1_13/U2  ( .A(
        \adder_0/operator_B_stage_1_13/n3 ), .ZN(\adder_0/G1[13] ) );
  AND2_X1 \adder_0/operator_B_stage_1_13/U1  ( .A1(\adder_0/P0[25] ), .A2(
        \adder_0/P0[26] ), .ZN(\adder_0/P1[13] ) );
  AOI21_X1 \adder_0/operator_B_stage_1_14/U3  ( .B1(\adder_0/G0[27] ), .B2(
        \adder_0/P0[28] ), .A(\adder_0/G0[28] ), .ZN(
        \adder_0/operator_B_stage_1_14/n3 ) );
  INV_X1 \adder_0/operator_B_stage_1_14/U2  ( .A(
        \adder_0/operator_B_stage_1_14/n3 ), .ZN(\adder_0/G1[14] ) );
  AND2_X1 \adder_0/operator_B_stage_1_14/U1  ( .A1(\adder_0/P0[27] ), .A2(
        \adder_0/P0[28] ), .ZN(\adder_0/P1[14] ) );
  AOI21_X1 \adder_0/operator_B_stage_1_15/U3  ( .B1(\adder_0/G0[29] ), .B2(
        \adder_0/P0[30] ), .A(\adder_0/G0[30] ), .ZN(
        \adder_0/operator_B_stage_1_15/n3 ) );
  INV_X1 \adder_0/operator_B_stage_1_15/U2  ( .A(
        \adder_0/operator_B_stage_1_15/n3 ), .ZN(\adder_0/G1[15] ) );
  AND2_X1 \adder_0/operator_B_stage_1_15/U1  ( .A1(\adder_0/P0[29] ), .A2(
        \adder_0/P0[30] ), .ZN(\adder_0/P1[15] ) );
  AOI21_X1 \adder_0/operator_C_stage_2_1/U2  ( .B1(\adder_0/P1[1] ), .B2(
        \adder_0/G1[0] ), .A(\adder_0/G1[1] ), .ZN(
        \adder_0/operator_C_stage_2_1/n3 ) );
  INV_X1 \adder_0/operator_C_stage_2_1/U1  ( .A(
        \adder_0/operator_C_stage_2_1/n3 ), .ZN(\adder_0/G2[1] ) );
  AOI21_X1 \adder_0/operator_B_stage_2_2/U3  ( .B1(\adder_0/G1[1] ), .B2(
        \adder_0/P1[2] ), .A(\adder_0/G1[2] ), .ZN(
        \adder_0/operator_B_stage_2_2/n3 ) );
  INV_X1 \adder_0/operator_B_stage_2_2/U2  ( .A(
        \adder_0/operator_B_stage_2_2/n3 ), .ZN(\adder_0/G2[2] ) );
  AND2_X1 \adder_0/operator_B_stage_2_2/U1  ( .A1(\adder_0/P1[1] ), .A2(
        \adder_0/P1[2] ), .ZN(\adder_0/P2[2] ) );
  AOI21_X1 \adder_0/operator_B_stage_2_3/U3  ( .B1(\adder_0/G1[2] ), .B2(
        \adder_0/P1[3] ), .A(\adder_0/G1[3] ), .ZN(
        \adder_0/operator_B_stage_2_3/n3 ) );
  INV_X1 \adder_0/operator_B_stage_2_3/U2  ( .A(
        \adder_0/operator_B_stage_2_3/n3 ), .ZN(\adder_0/G2[3] ) );
  AND2_X1 \adder_0/operator_B_stage_2_3/U1  ( .A1(\adder_0/P1[2] ), .A2(
        \adder_0/P1[3] ), .ZN(\adder_0/P2[3] ) );
  AOI21_X1 \adder_0/operator_B_stage_2_4/U3  ( .B1(\adder_0/G1[3] ), .B2(
        \adder_0/P1[4] ), .A(\adder_0/G1[4] ), .ZN(
        \adder_0/operator_B_stage_2_4/n3 ) );
  INV_X1 \adder_0/operator_B_stage_2_4/U2  ( .A(
        \adder_0/operator_B_stage_2_4/n3 ), .ZN(\adder_0/G2[4] ) );
  AND2_X1 \adder_0/operator_B_stage_2_4/U1  ( .A1(\adder_0/P1[3] ), .A2(
        \adder_0/P1[4] ), .ZN(\adder_0/P2[4] ) );
  AOI21_X1 \adder_0/operator_B_stage_2_5/U3  ( .B1(\adder_0/G1[4] ), .B2(
        \adder_0/P1[5] ), .A(\adder_0/G1[5] ), .ZN(
        \adder_0/operator_B_stage_2_5/n3 ) );
  INV_X1 \adder_0/operator_B_stage_2_5/U2  ( .A(
        \adder_0/operator_B_stage_2_5/n3 ), .ZN(\adder_0/G2[5] ) );
  AND2_X1 \adder_0/operator_B_stage_2_5/U1  ( .A1(\adder_0/P1[4] ), .A2(
        \adder_0/P1[5] ), .ZN(\adder_0/P2[5] ) );
  AOI21_X1 \adder_0/operator_B_stage_2_6/U3  ( .B1(\adder_0/G1[5] ), .B2(
        \adder_0/P1[6] ), .A(\adder_0/G1[6] ), .ZN(
        \adder_0/operator_B_stage_2_6/n3 ) );
  INV_X1 \adder_0/operator_B_stage_2_6/U2  ( .A(
        \adder_0/operator_B_stage_2_6/n3 ), .ZN(\adder_0/G2[6] ) );
  AND2_X1 \adder_0/operator_B_stage_2_6/U1  ( .A1(\adder_0/P1[5] ), .A2(
        \adder_0/P1[6] ), .ZN(\adder_0/P2[6] ) );
  AOI21_X1 \adder_0/operator_B_stage_2_7/U3  ( .B1(\adder_0/G1[6] ), .B2(
        \adder_0/P1[7] ), .A(\adder_0/G1[7] ), .ZN(
        \adder_0/operator_B_stage_2_7/n3 ) );
  INV_X1 \adder_0/operator_B_stage_2_7/U2  ( .A(
        \adder_0/operator_B_stage_2_7/n3 ), .ZN(\adder_0/G2[7] ) );
  AND2_X1 \adder_0/operator_B_stage_2_7/U1  ( .A1(\adder_0/P1[6] ), .A2(
        \adder_0/P1[7] ), .ZN(\adder_0/P2[7] ) );
  AOI21_X1 \adder_0/operator_B_stage_2_8/U3  ( .B1(\adder_0/G1[7] ), .B2(
        \adder_0/P1[8] ), .A(\adder_0/G1[8] ), .ZN(
        \adder_0/operator_B_stage_2_8/n3 ) );
  INV_X1 \adder_0/operator_B_stage_2_8/U2  ( .A(
        \adder_0/operator_B_stage_2_8/n3 ), .ZN(\adder_0/G2[8] ) );
  AND2_X1 \adder_0/operator_B_stage_2_8/U1  ( .A1(\adder_0/P1[7] ), .A2(
        \adder_0/P1[8] ), .ZN(\adder_0/P2[8] ) );
  AOI21_X1 \adder_0/operator_B_stage_2_9/U3  ( .B1(\adder_0/G1[8] ), .B2(
        \adder_0/P1[9] ), .A(\adder_0/G1[9] ), .ZN(
        \adder_0/operator_B_stage_2_9/n3 ) );
  INV_X1 \adder_0/operator_B_stage_2_9/U2  ( .A(
        \adder_0/operator_B_stage_2_9/n3 ), .ZN(\adder_0/G2[9] ) );
  AND2_X1 \adder_0/operator_B_stage_2_9/U1  ( .A1(\adder_0/P1[8] ), .A2(
        \adder_0/P1[9] ), .ZN(\adder_0/P2[9] ) );
  AOI21_X1 \adder_0/operator_B_stage_2_10/U3  ( .B1(\adder_0/G1[9] ), .B2(
        \adder_0/P1[10] ), .A(\adder_0/G1[10] ), .ZN(
        \adder_0/operator_B_stage_2_10/n3 ) );
  INV_X1 \adder_0/operator_B_stage_2_10/U2  ( .A(
        \adder_0/operator_B_stage_2_10/n3 ), .ZN(\adder_0/G2[10] ) );
  AND2_X1 \adder_0/operator_B_stage_2_10/U1  ( .A1(\adder_0/P1[9] ), .A2(
        \adder_0/P1[10] ), .ZN(\adder_0/P2[10] ) );
  AOI21_X1 \adder_0/operator_B_stage_2_11/U3  ( .B1(\adder_0/G1[10] ), .B2(
        \adder_0/P1[11] ), .A(\adder_0/G1[11] ), .ZN(
        \adder_0/operator_B_stage_2_11/n3 ) );
  INV_X1 \adder_0/operator_B_stage_2_11/U2  ( .A(
        \adder_0/operator_B_stage_2_11/n3 ), .ZN(\adder_0/G2[11] ) );
  AND2_X1 \adder_0/operator_B_stage_2_11/U1  ( .A1(\adder_0/P1[10] ), .A2(
        \adder_0/P1[11] ), .ZN(\adder_0/P2[11] ) );
  AOI21_X1 \adder_0/operator_B_stage_2_12/U3  ( .B1(\adder_0/G1[11] ), .B2(
        \adder_0/P1[12] ), .A(\adder_0/G1[12] ), .ZN(
        \adder_0/operator_B_stage_2_12/n3 ) );
  INV_X1 \adder_0/operator_B_stage_2_12/U2  ( .A(
        \adder_0/operator_B_stage_2_12/n3 ), .ZN(\adder_0/G2[12] ) );
  AND2_X1 \adder_0/operator_B_stage_2_12/U1  ( .A1(\adder_0/P1[11] ), .A2(
        \adder_0/P1[12] ), .ZN(\adder_0/P2[12] ) );
  AOI21_X1 \adder_0/operator_B_stage_2_13/U3  ( .B1(\adder_0/G1[12] ), .B2(
        \adder_0/P1[13] ), .A(\adder_0/G1[13] ), .ZN(
        \adder_0/operator_B_stage_2_13/n3 ) );
  INV_X1 \adder_0/operator_B_stage_2_13/U2  ( .A(
        \adder_0/operator_B_stage_2_13/n3 ), .ZN(\adder_0/G2[13] ) );
  AND2_X1 \adder_0/operator_B_stage_2_13/U1  ( .A1(\adder_0/P1[12] ), .A2(
        \adder_0/P1[13] ), .ZN(\adder_0/P2[13] ) );
  AOI21_X1 \adder_0/operator_B_stage_2_14/U3  ( .B1(\adder_0/G1[13] ), .B2(
        \adder_0/P1[14] ), .A(\adder_0/G1[14] ), .ZN(
        \adder_0/operator_B_stage_2_14/n3 ) );
  AND2_X1 \adder_0/operator_B_stage_2_14/U2  ( .A1(\adder_0/P1[13] ), .A2(
        \adder_0/P1[14] ), .ZN(\adder_0/P2[14] ) );
  INV_X1 \adder_0/operator_B_stage_2_14/U1  ( .A(
        \adder_0/operator_B_stage_2_14/n3 ), .ZN(\adder_0/G2[14] ) );
  AOI21_X1 \adder_0/operator_B_stage_2_15/U3  ( .B1(\adder_0/G1[14] ), .B2(
        \adder_0/P1[15] ), .A(\adder_0/G1[15] ), .ZN(
        \adder_0/operator_B_stage_2_15/n3 ) );
  INV_X1 \adder_0/operator_B_stage_2_15/U2  ( .A(
        \adder_0/operator_B_stage_2_15/n3 ), .ZN(\adder_0/G2[15] ) );
  AND2_X1 \adder_0/operator_B_stage_2_15/U1  ( .A1(\adder_0/P1[14] ), .A2(
        \adder_0/P1[15] ), .ZN(\adder_0/P2[15] ) );
  AOI21_X1 \adder_0/operator_C_stage_3_2/U2  ( .B1(\adder_0/P2[2] ), .B2(
        \adder_0/G1[0] ), .A(\adder_0/G2[2] ), .ZN(
        \adder_0/operator_C_stage_3_2/n3 ) );
  INV_X1 \adder_0/operator_C_stage_3_2/U1  ( .A(
        \adder_0/operator_C_stage_3_2/n3 ), .ZN(\adder_0/G3[2] ) );
  AOI21_X1 \adder_0/operator_C_stage_3_3/U2  ( .B1(\adder_0/P2[3] ), .B2(
        \adder_0/G2[1] ), .A(\adder_0/G2[3] ), .ZN(
        \adder_0/operator_C_stage_3_3/n3 ) );
  INV_X1 \adder_0/operator_C_stage_3_3/U1  ( .A(
        \adder_0/operator_C_stage_3_3/n3 ), .ZN(\adder_0/G3[3] ) );
  AOI21_X1 \adder_0/operator_B_stage_3_4/U3  ( .B1(\adder_0/G2[2] ), .B2(
        \adder_0/P2[4] ), .A(\adder_0/G2[4] ), .ZN(
        \adder_0/operator_B_stage_3_4/n3 ) );
  INV_X1 \adder_0/operator_B_stage_3_4/U2  ( .A(
        \adder_0/operator_B_stage_3_4/n3 ), .ZN(\adder_0/G3[4] ) );
  AND2_X1 \adder_0/operator_B_stage_3_4/U1  ( .A1(\adder_0/P2[2] ), .A2(
        \adder_0/P2[4] ), .ZN(\adder_0/P3[4] ) );
  AOI21_X1 \adder_0/operator_B_stage_3_5/U3  ( .B1(\adder_0/G2[3] ), .B2(
        \adder_0/P2[5] ), .A(\adder_0/G2[5] ), .ZN(
        \adder_0/operator_B_stage_3_5/n3 ) );
  INV_X1 \adder_0/operator_B_stage_3_5/U2  ( .A(
        \adder_0/operator_B_stage_3_5/n3 ), .ZN(\adder_0/G3[5] ) );
  AND2_X1 \adder_0/operator_B_stage_3_5/U1  ( .A1(\adder_0/P2[3] ), .A2(
        \adder_0/P2[5] ), .ZN(\adder_0/P3[5] ) );
  AOI21_X1 \adder_0/operator_B_stage_3_6/U3  ( .B1(\adder_0/G2[4] ), .B2(
        \adder_0/P2[6] ), .A(\adder_0/G2[6] ), .ZN(
        \adder_0/operator_B_stage_3_6/n3 ) );
  INV_X1 \adder_0/operator_B_stage_3_6/U2  ( .A(
        \adder_0/operator_B_stage_3_6/n3 ), .ZN(\adder_0/G3[6] ) );
  AND2_X1 \adder_0/operator_B_stage_3_6/U1  ( .A1(\adder_0/P2[4] ), .A2(
        \adder_0/P2[6] ), .ZN(\adder_0/P3[6] ) );
  AOI21_X1 \adder_0/operator_B_stage_3_7/U3  ( .B1(\adder_0/G2[5] ), .B2(
        \adder_0/P2[7] ), .A(\adder_0/G2[7] ), .ZN(
        \adder_0/operator_B_stage_3_7/n3 ) );
  INV_X1 \adder_0/operator_B_stage_3_7/U2  ( .A(
        \adder_0/operator_B_stage_3_7/n3 ), .ZN(\adder_0/G3[7] ) );
  AND2_X1 \adder_0/operator_B_stage_3_7/U1  ( .A1(\adder_0/P2[5] ), .A2(
        \adder_0/P2[7] ), .ZN(\adder_0/P3[7] ) );
  AOI21_X1 \adder_0/operator_B_stage_3_8/U3  ( .B1(\adder_0/G2[6] ), .B2(
        \adder_0/P2[8] ), .A(\adder_0/G2[8] ), .ZN(
        \adder_0/operator_B_stage_3_8/n3 ) );
  INV_X1 \adder_0/operator_B_stage_3_8/U2  ( .A(
        \adder_0/operator_B_stage_3_8/n3 ), .ZN(\adder_0/G3[8] ) );
  AND2_X1 \adder_0/operator_B_stage_3_8/U1  ( .A1(\adder_0/P2[6] ), .A2(
        \adder_0/P2[8] ), .ZN(\adder_0/P3[8] ) );
  AOI21_X1 \adder_0/operator_B_stage_3_9/U3  ( .B1(\adder_0/G2[7] ), .B2(
        \adder_0/P2[9] ), .A(\adder_0/G2[9] ), .ZN(
        \adder_0/operator_B_stage_3_9/n3 ) );
  INV_X1 \adder_0/operator_B_stage_3_9/U2  ( .A(
        \adder_0/operator_B_stage_3_9/n3 ), .ZN(\adder_0/G3[9] ) );
  AND2_X1 \adder_0/operator_B_stage_3_9/U1  ( .A1(\adder_0/P2[7] ), .A2(
        \adder_0/P2[9] ), .ZN(\adder_0/P3[9] ) );
  AOI21_X1 \adder_0/operator_B_stage_3_10/U3  ( .B1(\adder_0/G2[8] ), .B2(
        \adder_0/P2[10] ), .A(\adder_0/G2[10] ), .ZN(
        \adder_0/operator_B_stage_3_10/n3 ) );
  INV_X1 \adder_0/operator_B_stage_3_10/U2  ( .A(
        \adder_0/operator_B_stage_3_10/n3 ), .ZN(\adder_0/G3[10] ) );
  AND2_X1 \adder_0/operator_B_stage_3_10/U1  ( .A1(\adder_0/P2[8] ), .A2(
        \adder_0/P2[10] ), .ZN(\adder_0/P3[10] ) );
  AOI21_X1 \adder_0/operator_B_stage_3_11/U3  ( .B1(\adder_0/G2[9] ), .B2(
        \adder_0/P2[11] ), .A(\adder_0/G2[11] ), .ZN(
        \adder_0/operator_B_stage_3_11/n3 ) );
  INV_X1 \adder_0/operator_B_stage_3_11/U2  ( .A(
        \adder_0/operator_B_stage_3_11/n3 ), .ZN(\adder_0/G3[11] ) );
  AND2_X1 \adder_0/operator_B_stage_3_11/U1  ( .A1(\adder_0/P2[9] ), .A2(
        \adder_0/P2[11] ), .ZN(\adder_0/P3[11] ) );
  AOI21_X1 \adder_0/operator_B_stage_3_12/U3  ( .B1(\adder_0/G2[10] ), .B2(
        \adder_0/P2[12] ), .A(\adder_0/G2[12] ), .ZN(
        \adder_0/operator_B_stage_3_12/n3 ) );
  INV_X1 \adder_0/operator_B_stage_3_12/U2  ( .A(
        \adder_0/operator_B_stage_3_12/n3 ), .ZN(\adder_0/G3[12] ) );
  AND2_X1 \adder_0/operator_B_stage_3_12/U1  ( .A1(\adder_0/P2[10] ), .A2(
        \adder_0/P2[12] ), .ZN(\adder_0/P3[12] ) );
  AOI21_X1 \adder_0/operator_B_stage_3_13/U3  ( .B1(\adder_0/G2[11] ), .B2(
        \adder_0/P2[13] ), .A(\adder_0/G2[13] ), .ZN(
        \adder_0/operator_B_stage_3_13/n3 ) );
  INV_X1 \adder_0/operator_B_stage_3_13/U2  ( .A(
        \adder_0/operator_B_stage_3_13/n3 ), .ZN(\adder_0/G3[13] ) );
  AND2_X1 \adder_0/operator_B_stage_3_13/U1  ( .A1(\adder_0/P2[11] ), .A2(
        \adder_0/P2[13] ), .ZN(\adder_0/P3[13] ) );
  AOI21_X1 \adder_0/operator_B_stage_3_14/U3  ( .B1(\adder_0/G2[12] ), .B2(
        \adder_0/P2[14] ), .A(\adder_0/G2[14] ), .ZN(
        \adder_0/operator_B_stage_3_14/n3 ) );
  INV_X1 \adder_0/operator_B_stage_3_14/U2  ( .A(
        \adder_0/operator_B_stage_3_14/n3 ), .ZN(\adder_0/G3[14] ) );
  AND2_X1 \adder_0/operator_B_stage_3_14/U1  ( .A1(\adder_0/P2[12] ), .A2(
        \adder_0/P2[14] ), .ZN(\adder_0/P3[14] ) );
  AOI21_X1 \adder_0/operator_B_stage_3_15/U3  ( .B1(\adder_0/G2[13] ), .B2(
        \adder_0/P2[15] ), .A(\adder_0/G2[15] ), .ZN(
        \adder_0/operator_B_stage_3_15/n3 ) );
  INV_X1 \adder_0/operator_B_stage_3_15/U2  ( .A(
        \adder_0/operator_B_stage_3_15/n3 ), .ZN(\adder_0/G3[15] ) );
  AND2_X1 \adder_0/operator_B_stage_3_15/U1  ( .A1(\adder_0/P2[13] ), .A2(
        \adder_0/P2[15] ), .ZN(\adder_0/P3[15] ) );
  AOI21_X1 \adder_0/operator_C_stage_4_4/U2  ( .B1(\adder_0/P3[4] ), .B2(
        \adder_0/G1[0] ), .A(\adder_0/G3[4] ), .ZN(
        \adder_0/operator_C_stage_4_4/n3 ) );
  INV_X1 \adder_0/operator_C_stage_4_4/U1  ( .A(
        \adder_0/operator_C_stage_4_4/n3 ), .ZN(\adder_0/G4[4] ) );
  AOI21_X1 \adder_0/operator_C_stage_4_5/U2  ( .B1(\adder_0/P3[5] ), .B2(
        \adder_0/G2[1] ), .A(\adder_0/G3[5] ), .ZN(
        \adder_0/operator_C_stage_4_5/n3 ) );
  INV_X1 \adder_0/operator_C_stage_4_5/U1  ( .A(
        \adder_0/operator_C_stage_4_5/n3 ), .ZN(\adder_0/G4[5] ) );
  AOI21_X1 \adder_0/operator_C_stage_4_6/U2  ( .B1(\adder_0/P3[6] ), .B2(
        \adder_0/G3[2] ), .A(\adder_0/G3[6] ), .ZN(
        \adder_0/operator_C_stage_4_6/n3 ) );
  INV_X1 \adder_0/operator_C_stage_4_6/U1  ( .A(
        \adder_0/operator_C_stage_4_6/n3 ), .ZN(\adder_0/G4[6] ) );
  AOI21_X1 \adder_0/operator_C_stage_4_7/U2  ( .B1(\adder_0/P3[7] ), .B2(
        \adder_0/G3[3] ), .A(\adder_0/G3[7] ), .ZN(
        \adder_0/operator_C_stage_4_7/n3 ) );
  INV_X1 \adder_0/operator_C_stage_4_7/U1  ( .A(
        \adder_0/operator_C_stage_4_7/n3 ), .ZN(\adder_0/G4[7] ) );
  INV_X1 \adder_0/operator_B_stage_4_8/U3  ( .A(
        \adder_0/operator_B_stage_4_8/n3 ), .ZN(\adder_0/G4[8] ) );
  AND2_X1 \adder_0/operator_B_stage_4_8/U2  ( .A1(\adder_0/P3[4] ), .A2(
        \adder_0/P3[8] ), .ZN(\adder_0/P4 [8]) );
  AOI21_X1 \adder_0/operator_B_stage_4_8/U1  ( .B1(\adder_0/G3[4] ), .B2(
        \adder_0/P3[8] ), .A(\adder_0/G3[8] ), .ZN(
        \adder_0/operator_B_stage_4_8/n3 ) );
  INV_X1 \adder_0/operator_B_stage_4_9/U3  ( .A(
        \adder_0/operator_B_stage_4_9/n3 ), .ZN(\adder_0/G4[9] ) );
  AND2_X1 \adder_0/operator_B_stage_4_9/U2  ( .A1(\adder_0/P3[5] ), .A2(
        \adder_0/P3[9] ), .ZN(\adder_0/P4 [9]) );
  AOI21_X1 \adder_0/operator_B_stage_4_9/U1  ( .B1(\adder_0/G3[5] ), .B2(
        \adder_0/P3[9] ), .A(\adder_0/G3[9] ), .ZN(
        \adder_0/operator_B_stage_4_9/n3 ) );
  INV_X1 \adder_0/operator_B_stage_4_10/U3  ( .A(
        \adder_0/operator_B_stage_4_10/n3 ), .ZN(\adder_0/G4[10] ) );
  AND2_X1 \adder_0/operator_B_stage_4_10/U2  ( .A1(\adder_0/P3[6] ), .A2(
        \adder_0/P3[10] ), .ZN(\adder_0/P4 [10]) );
  AOI21_X1 \adder_0/operator_B_stage_4_10/U1  ( .B1(\adder_0/G3[6] ), .B2(
        \adder_0/P3[10] ), .A(\adder_0/G3[10] ), .ZN(
        \adder_0/operator_B_stage_4_10/n3 ) );
  INV_X1 \adder_0/operator_B_stage_4_11/U3  ( .A(
        \adder_0/operator_B_stage_4_11/n3 ), .ZN(\adder_0/G4[11] ) );
  AND2_X1 \adder_0/operator_B_stage_4_11/U2  ( .A1(\adder_0/P3[7] ), .A2(
        \adder_0/P3[11] ), .ZN(\adder_0/P4 [11]) );
  AOI21_X1 \adder_0/operator_B_stage_4_11/U1  ( .B1(\adder_0/G3[7] ), .B2(
        \adder_0/P3[11] ), .A(\adder_0/G3[11] ), .ZN(
        \adder_0/operator_B_stage_4_11/n3 ) );
  INV_X1 \adder_0/operator_B_stage_4_12/U3  ( .A(
        \adder_0/operator_B_stage_4_12/n3 ), .ZN(\adder_0/G4[12] ) );
  AND2_X1 \adder_0/operator_B_stage_4_12/U2  ( .A1(\adder_0/P3[8] ), .A2(
        \adder_0/P3[12] ), .ZN(\adder_0/P4 [12]) );
  AOI21_X1 \adder_0/operator_B_stage_4_12/U1  ( .B1(\adder_0/G3[8] ), .B2(
        \adder_0/P3[12] ), .A(\adder_0/G3[12] ), .ZN(
        \adder_0/operator_B_stage_4_12/n3 ) );
  AOI21_X1 \adder_0/operator_B_stage_4_13/U3  ( .B1(\adder_0/G3[9] ), .B2(
        \adder_0/P3[13] ), .A(\adder_0/G3[13] ), .ZN(
        \adder_0/operator_B_stage_4_13/n3 ) );
  INV_X1 \adder_0/operator_B_stage_4_13/U2  ( .A(
        \adder_0/operator_B_stage_4_13/n3 ), .ZN(\adder_0/G4[13] ) );
  AND2_X1 \adder_0/operator_B_stage_4_13/U1  ( .A1(\adder_0/P3[9] ), .A2(
        \adder_0/P3[13] ), .ZN(\adder_0/P4 [13]) );
  AOI21_X1 \adder_0/operator_B_stage_4_14/U3  ( .B1(\adder_0/G3[10] ), .B2(
        \adder_0/P3[14] ), .A(\adder_0/G3[14] ), .ZN(
        \adder_0/operator_B_stage_4_14/n3 ) );
  INV_X1 \adder_0/operator_B_stage_4_14/U2  ( .A(
        \adder_0/operator_B_stage_4_14/n3 ), .ZN(\adder_0/G4[14] ) );
  AND2_X1 \adder_0/operator_B_stage_4_14/U1  ( .A1(\adder_0/P3[10] ), .A2(
        \adder_0/P3[14] ), .ZN(\adder_0/P4 [14]) );
  AOI21_X1 \adder_0/operator_B_stage_4_15/U3  ( .B1(\adder_0/G3[11] ), .B2(
        \adder_0/P3[15] ), .A(\adder_0/G3[15] ), .ZN(
        \adder_0/operator_B_stage_4_15/n3 ) );
  INV_X1 \adder_0/operator_B_stage_4_15/U2  ( .A(
        \adder_0/operator_B_stage_4_15/n3 ), .ZN(\adder_0/G4[15] ) );
  AND2_X1 \adder_0/operator_B_stage_4_15/U1  ( .A1(\adder_0/P3[11] ), .A2(
        \adder_0/P3[15] ), .ZN(\adder_0/P4 [15]) );
  AOI21_X1 \adder_0/operator_C_stage_5_8/U2  ( .B1(\adder_0/P4 [8]), .B2(
        \adder_0/G1[0] ), .A(\adder_0/G4[8] ), .ZN(
        \adder_0/operator_C_stage_5_8/n3 ) );
  INV_X1 \adder_0/operator_C_stage_5_8/U1  ( .A(
        \adder_0/operator_C_stage_5_8/n3 ), .ZN(\adder_0/G5[8] ) );
  AOI21_X1 \adder_0/operator_C_stage_5_9/U2  ( .B1(\adder_0/P4 [9]), .B2(
        \adder_0/G2[1] ), .A(\adder_0/G4[9] ), .ZN(
        \adder_0/operator_C_stage_5_9/n3 ) );
  INV_X1 \adder_0/operator_C_stage_5_9/U1  ( .A(
        \adder_0/operator_C_stage_5_9/n3 ), .ZN(\adder_0/G5[9] ) );
  AOI21_X1 \adder_0/operator_C_stage_5_10/U2  ( .B1(\adder_0/P4 [10]), .B2(
        \adder_0/G3[2] ), .A(\adder_0/G4[10] ), .ZN(
        \adder_0/operator_C_stage_5_10/n3 ) );
  INV_X1 \adder_0/operator_C_stage_5_10/U1  ( .A(
        \adder_0/operator_C_stage_5_10/n3 ), .ZN(\adder_0/G5[10] ) );
  AOI21_X1 \adder_0/operator_C_stage_5_11/U2  ( .B1(\adder_0/P4 [11]), .B2(
        \adder_0/G3[3] ), .A(\adder_0/G4[11] ), .ZN(
        \adder_0/operator_C_stage_5_11/n3 ) );
  INV_X1 \adder_0/operator_C_stage_5_11/U1  ( .A(
        \adder_0/operator_C_stage_5_11/n3 ), .ZN(\adder_0/G5[11] ) );
  AOI21_X1 \adder_0/operator_C_stage_5_12/U2  ( .B1(\adder_0/P4 [12]), .B2(
        \adder_0/G4[4] ), .A(\adder_0/G4[12] ), .ZN(
        \adder_0/operator_C_stage_5_12/n3 ) );
  INV_X1 \adder_0/operator_C_stage_5_12/U1  ( .A(
        \adder_0/operator_C_stage_5_12/n3 ), .ZN(\adder_0/G5[12] ) );
  AOI21_X1 \adder_0/operator_C_stage_5_13/U2  ( .B1(\adder_0/P4 [13]), .B2(
        \adder_0/G4[5] ), .A(\adder_0/G4[13] ), .ZN(
        \adder_0/operator_C_stage_5_13/n3 ) );
  INV_X1 \adder_0/operator_C_stage_5_13/U1  ( .A(
        \adder_0/operator_C_stage_5_13/n3 ), .ZN(\adder_0/G5[13] ) );
  AOI21_X1 \adder_0/operator_C_stage_5_14/U2  ( .B1(\adder_0/P4 [14]), .B2(
        \adder_0/G4[6] ), .A(\adder_0/G4[14] ), .ZN(
        \adder_0/operator_C_stage_5_14/n3 ) );
  INV_X1 \adder_0/operator_C_stage_5_14/U1  ( .A(
        \adder_0/operator_C_stage_5_14/n3 ), .ZN(\adder_0/G5[14] ) );
  AOI21_X1 \adder_0/operator_C_stage_5_15/U2  ( .B1(\adder_0/P4 [15]), .B2(
        \adder_0/G4[7] ), .A(\adder_0/G4[15] ), .ZN(
        \adder_0/operator_C_stage_5_15/n3 ) );
  INV_X1 \adder_0/operator_C_stage_5_15/U1  ( .A(
        \adder_0/operator_C_stage_5_15/n3 ), .ZN(\adder_0/G5[15] ) );
  AOI21_X1 \adder_0/operator_C_stage_6_0/U2  ( .B1(\adder_0/P0[1] ), .B2(
        \adder_0/G1[0] ), .A(\adder_0/G0[1] ), .ZN(
        \adder_0/operator_C_stage_6_0/n3 ) );
  INV_X1 \adder_0/operator_C_stage_6_0/U1  ( .A(
        \adder_0/operator_C_stage_6_0/n3 ), .ZN(\adder_0/G6_1 ) );
  AOI21_X1 \adder_0/operator_C_stage_6_1/U2  ( .B1(\adder_0/P0[3] ), .B2(
        \adder_0/G2[1] ), .A(\adder_0/G0[3] ), .ZN(
        \adder_0/operator_C_stage_6_1/n3 ) );
  INV_X1 \adder_0/operator_C_stage_6_1/U1  ( .A(
        \adder_0/operator_C_stage_6_1/n3 ), .ZN(\adder_0/G6_3 ) );
  AOI21_X1 \adder_0/operator_C_stage_6_2/U2  ( .B1(\adder_0/P0[5] ), .B2(
        \adder_0/G3[2] ), .A(\adder_0/G0[5] ), .ZN(
        \adder_0/operator_C_stage_6_2/n3 ) );
  INV_X1 \adder_0/operator_C_stage_6_2/U1  ( .A(
        \adder_0/operator_C_stage_6_2/n3 ), .ZN(\adder_0/G6_5 ) );
  AOI21_X1 \adder_0/operator_C_stage_6_3/U2  ( .B1(\adder_0/P0[7] ), .B2(
        \adder_0/G3[3] ), .A(\adder_0/G0[7] ), .ZN(
        \adder_0/operator_C_stage_6_3/n3 ) );
  INV_X1 \adder_0/operator_C_stage_6_3/U1  ( .A(
        \adder_0/operator_C_stage_6_3/n3 ), .ZN(\adder_0/G6_7 ) );
  AOI21_X1 \adder_0/operator_C_stage_6_4/U2  ( .B1(\adder_0/P0[9] ), .B2(
        \adder_0/G4[4] ), .A(\adder_0/G0[9] ), .ZN(
        \adder_0/operator_C_stage_6_4/n3 ) );
  INV_X1 \adder_0/operator_C_stage_6_4/U1  ( .A(
        \adder_0/operator_C_stage_6_4/n3 ), .ZN(\adder_0/G6_9 ) );
  AOI21_X1 \adder_0/operator_C_stage_6_5/U2  ( .B1(\adder_0/P0[11] ), .B2(
        \adder_0/G4[5] ), .A(\adder_0/G0[11] ), .ZN(
        \adder_0/operator_C_stage_6_5/n3 ) );
  INV_X1 \adder_0/operator_C_stage_6_5/U1  ( .A(
        \adder_0/operator_C_stage_6_5/n3 ), .ZN(\adder_0/G6_11 ) );
  AOI21_X1 \adder_0/operator_C_stage_6_6/U2  ( .B1(\adder_0/P0[13] ), .B2(
        \adder_0/G4[6] ), .A(\adder_0/G0[13] ), .ZN(
        \adder_0/operator_C_stage_6_6/n3 ) );
  INV_X1 \adder_0/operator_C_stage_6_6/U1  ( .A(
        \adder_0/operator_C_stage_6_6/n3 ), .ZN(\adder_0/G6_13 ) );
  AOI21_X1 \adder_0/operator_C_stage_6_7/U2  ( .B1(\adder_0/P0[15] ), .B2(
        \adder_0/G4[7] ), .A(\adder_0/G0[15] ), .ZN(
        \adder_0/operator_C_stage_6_7/n3 ) );
  INV_X1 \adder_0/operator_C_stage_6_7/U1  ( .A(
        \adder_0/operator_C_stage_6_7/n3 ), .ZN(\adder_0/G6_15 ) );
  AOI21_X1 \adder_0/operator_C_stage_6_8/U2  ( .B1(\adder_0/P0[17] ), .B2(
        \adder_0/G5[8] ), .A(\adder_0/G0[17] ), .ZN(
        \adder_0/operator_C_stage_6_8/n3 ) );
  INV_X1 \adder_0/operator_C_stage_6_8/U1  ( .A(
        \adder_0/operator_C_stage_6_8/n3 ), .ZN(\adder_0/G6_17 ) );
  AOI21_X1 \adder_0/operator_C_stage_6_9/U2  ( .B1(\adder_0/P0[19] ), .B2(
        \adder_0/G5[9] ), .A(\adder_0/G0[19] ), .ZN(
        \adder_0/operator_C_stage_6_9/n3 ) );
  INV_X1 \adder_0/operator_C_stage_6_9/U1  ( .A(
        \adder_0/operator_C_stage_6_9/n3 ), .ZN(\adder_0/G6_19 ) );
  AOI21_X1 \adder_0/operator_C_stage_6_10/U2  ( .B1(\adder_0/P0[21] ), .B2(
        \adder_0/G5[10] ), .A(\adder_0/G0[21] ), .ZN(
        \adder_0/operator_C_stage_6_10/n3 ) );
  INV_X1 \adder_0/operator_C_stage_6_10/U1  ( .A(
        \adder_0/operator_C_stage_6_10/n3 ), .ZN(\adder_0/G6_21 ) );
  AOI21_X1 \adder_0/operator_C_stage_6_11/U2  ( .B1(\adder_0/P0[23] ), .B2(
        \adder_0/G5[11] ), .A(\adder_0/G0[23] ), .ZN(
        \adder_0/operator_C_stage_6_11/n3 ) );
  INV_X1 \adder_0/operator_C_stage_6_11/U1  ( .A(
        \adder_0/operator_C_stage_6_11/n3 ), .ZN(\adder_0/G6_23 ) );
  AOI21_X1 \adder_0/operator_C_stage_6_12/U2  ( .B1(\adder_0/P0[25] ), .B2(
        \adder_0/G5[12] ), .A(\adder_0/G0[25] ), .ZN(
        \adder_0/operator_C_stage_6_12/n3 ) );
  INV_X1 \adder_0/operator_C_stage_6_12/U1  ( .A(
        \adder_0/operator_C_stage_6_12/n3 ), .ZN(\adder_0/G6_25 ) );
  AOI21_X1 \adder_0/operator_C_stage_6_13/U2  ( .B1(\adder_0/P0[27] ), .B2(
        \adder_0/G5[13] ), .A(\adder_0/G0[27] ), .ZN(
        \adder_0/operator_C_stage_6_13/n3 ) );
  INV_X1 \adder_0/operator_C_stage_6_13/U1  ( .A(
        \adder_0/operator_C_stage_6_13/n3 ), .ZN(\adder_0/G6_27 ) );
  AOI21_X1 \adder_0/operator_C_stage_6_14/U2  ( .B1(\adder_0/P0[29] ), .B2(
        \adder_0/G5[14] ), .A(\adder_0/G0[29] ), .ZN(
        \adder_0/operator_C_stage_6_14/n3 ) );
  INV_X1 \adder_0/operator_C_stage_6_14/U1  ( .A(
        \adder_0/operator_C_stage_6_14/n3 ), .ZN(\adder_0/G6_29_ ) );
  AOI21_X1 \adder_0/operator_C_stage_6_15/U2  ( .B1(\adder_0/P0[31] ), .B2(
        \adder_0/G5[15] ), .A(\adder_0/G0[31] ), .ZN(
        \adder_0/operator_C_stage_6_15/n3 ) );
  INV_X1 \adder_0/operator_C_stage_6_15/U1  ( .A(
        \adder_0/operator_C_stage_6_15/n3 ), .ZN(\adder_0/o_c ) );
  XOR2_X1 \adder_1/U32  ( .A(n2983), .B(\adder_1/P0[0] ), .Z(sum_ct[0]) );
  XOR2_X1 \adder_1/U31  ( .A(\adder_1/P0[10] ), .B(\adder_1/G6_9 ), .Z(
        SYNOPSYS_UNCONNECTED_23) );
  XOR2_X1 \adder_1/U30  ( .A(\adder_1/P0[11] ), .B(\adder_1/G4[5] ), .Z(
        SYNOPSYS_UNCONNECTED_22) );
  XOR2_X1 \adder_1/U29  ( .A(\adder_1/P0[12] ), .B(\adder_1/G6_11 ), .Z(
        SYNOPSYS_UNCONNECTED_21) );
  XOR2_X1 \adder_1/U28  ( .A(\adder_1/P0[13] ), .B(\adder_1/G4[6] ), .Z(
        SYNOPSYS_UNCONNECTED_20) );
  XOR2_X1 \adder_1/U27  ( .A(\adder_1/P0[14] ), .B(\adder_1/G6_13 ), .Z(
        SYNOPSYS_UNCONNECTED_19) );
  XOR2_X1 \adder_1/U26  ( .A(\adder_1/P0[15] ), .B(\adder_1/G4[7] ), .Z(
        SYNOPSYS_UNCONNECTED_18) );
  XOR2_X1 \adder_1/U25  ( .A(\adder_1/P0[16] ), .B(\adder_1/G6_15 ), .Z(
        SYNOPSYS_UNCONNECTED_17) );
  XOR2_X1 \adder_1/U24  ( .A(\adder_1/P0[17] ), .B(\adder_1/G5[8] ), .Z(
        SYNOPSYS_UNCONNECTED_16) );
  XOR2_X1 \adder_1/U23  ( .A(\adder_1/P0[18] ), .B(\adder_1/G6_17 ), .Z(
        SYNOPSYS_UNCONNECTED_15) );
  XOR2_X1 \adder_1/U22  ( .A(\adder_1/P0[19] ), .B(\adder_1/G5[9] ), .Z(
        SYNOPSYS_UNCONNECTED_14) );
  XOR2_X1 \adder_1/U21  ( .A(\adder_1/P0[1] ), .B(\adder_1/G1[0] ), .Z(
        sum_ct[1]) );
  XOR2_X1 \adder_1/U20  ( .A(\adder_1/P0[20] ), .B(\adder_1/G6_19 ), .Z(
        SYNOPSYS_UNCONNECTED_13) );
  XOR2_X1 \adder_1/U19  ( .A(\adder_1/P0[21] ), .B(\adder_1/G5[10] ), .Z(
        SYNOPSYS_UNCONNECTED_12) );
  XOR2_X1 \adder_1/U18  ( .A(\adder_1/P0[22] ), .B(\adder_1/G6_21 ), .Z(
        SYNOPSYS_UNCONNECTED_11) );
  XOR2_X1 \adder_1/U17  ( .A(\adder_1/P0[23] ), .B(\adder_1/G5[11] ), .Z(
        SYNOPSYS_UNCONNECTED_10) );
  XOR2_X1 \adder_1/U16  ( .A(\adder_1/P0[24] ), .B(\adder_1/G6_23 ), .Z(
        SYNOPSYS_UNCONNECTED_9) );
  XOR2_X1 \adder_1/U15  ( .A(\adder_1/P0[25] ), .B(\adder_1/G5[12] ), .Z(
        SYNOPSYS_UNCONNECTED_8) );
  XOR2_X1 \adder_1/U14  ( .A(\adder_1/P0[26] ), .B(\adder_1/G6_25 ), .Z(
        SYNOPSYS_UNCONNECTED_7) );
  XOR2_X1 \adder_1/U13  ( .A(\adder_1/P0[27] ), .B(\adder_1/G5[13] ), .Z(
        SYNOPSYS_UNCONNECTED_6) );
  XOR2_X1 \adder_1/U12  ( .A(\adder_1/P0[28] ), .B(\adder_1/G6_27 ), .Z(
        SYNOPSYS_UNCONNECTED_5) );
  XOR2_X1 \adder_1/U11  ( .A(\adder_1/P0[29] ), .B(\adder_1/G5[14] ), .Z(
        SYNOPSYS_UNCONNECTED_4) );
  XOR2_X1 \adder_1/U10  ( .A(\adder_1/P0[2] ), .B(\adder_1/G6_1 ), .Z(
        sum_ct[2]) );
  XOR2_X1 \adder_1/U9  ( .A(\adder_1/P0[30] ), .B(\adder_1/G6_29_ ), .Z(
        SYNOPSYS_UNCONNECTED_3) );
  XOR2_X1 \adder_1/U8  ( .A(\adder_1/P0[31] ), .B(\adder_1/G5[15] ), .Z(
        SYNOPSYS_UNCONNECTED_2) );
  XOR2_X1 \adder_1/U7  ( .A(\adder_1/P0[3] ), .B(\adder_1/G2[1] ), .Z(
        sum_ct[3]) );
  XOR2_X1 \adder_1/U6  ( .A(\adder_1/P0[4] ), .B(\adder_1/G6_3 ), .Z(sum_ct[4]) );
  XOR2_X1 \adder_1/U5  ( .A(\adder_1/P0[5] ), .B(\adder_1/G3[2] ), .Z(
        sum_ct[5]) );
  XOR2_X1 \adder_1/U4  ( .A(\adder_1/P0[6] ), .B(\adder_1/G6_5 ), .Z(
        SYNOPSYS_UNCONNECTED_27) );
  XOR2_X1 \adder_1/U3  ( .A(\adder_1/P0[7] ), .B(\adder_1/G3[3] ), .Z(
        SYNOPSYS_UNCONNECTED_26) );
  XOR2_X1 \adder_1/U2  ( .A(\adder_1/P0[8] ), .B(\adder_1/G6_7 ), .Z(
        SYNOPSYS_UNCONNECTED_25) );
  XOR2_X1 \adder_1/U1  ( .A(\adder_1/P0[9] ), .B(\adder_1/G4[4] ), .Z(
        SYNOPSYS_UNCONNECTED_24) );
  AND2_X1 \adder_1/operator_A_0/U1  ( .A1(n_1_net__0_), .A2(ct[0]), .ZN(
        \adder_1/G0[0] ) );
  XOR2_X1 \adder_1/operator_A_0/U2  ( .A(n_1_net__0_), .B(ct[0]), .Z(
        \adder_1/P0[0] ) );
  AND2_X1 \adder_1/operator_A_1/U1  ( .A1(n_1_net__1_), .A2(ct[1]), .ZN(
        \adder_1/G0[1] ) );
  XOR2_X1 \adder_1/operator_A_1/U2  ( .A(n_1_net__1_), .B(ct[1]), .Z(
        \adder_1/P0[1] ) );
  AND2_X1 \adder_1/operator_A_2/U1  ( .A1(n_1_net__2_), .A2(ct[2]), .ZN(
        \adder_1/G0[2] ) );
  XOR2_X1 \adder_1/operator_A_2/U2  ( .A(n_1_net__2_), .B(ct[2]), .Z(
        \adder_1/P0[2] ) );
  AND2_X1 \adder_1/operator_A_3/U1  ( .A1(n_1_net__3_), .A2(ct[3]), .ZN(
        \adder_1/G0[3] ) );
  XOR2_X1 \adder_1/operator_A_3/U2  ( .A(n_1_net__3_), .B(ct[3]), .Z(
        \adder_1/P0[3] ) );
  AND2_X1 \adder_1/operator_A_4/U1  ( .A1(n2983), .A2(ct[4]), .ZN(
        \adder_1/G0[4] ) );
  XOR2_X1 \adder_1/operator_A_4/U2  ( .A(n2983), .B(ct[4]), .Z(\adder_1/P0[4] ) );
  AND2_X1 \adder_1/operator_A_5/U1  ( .A1(n2983), .A2(ct[5]), .ZN(
        \adder_1/G0[5] ) );
  XOR2_X1 \adder_1/operator_A_5/U2  ( .A(n2983), .B(ct[5]), .Z(\adder_1/P0[5] ) );
  AND2_X1 \adder_1/operator_A_6/U1  ( .A1(n2983), .A2(1'b0), .ZN(
        \adder_1/G0[6] ) );
  XOR2_X1 \adder_1/operator_A_6/U2  ( .A(n2983), .B(1'b0), .Z(\adder_1/P0[6] )
         );
  AND2_X1 \adder_1/operator_A_7/U1  ( .A1(n2983), .A2(1'b0), .ZN(
        \adder_1/G0[7] ) );
  XOR2_X1 \adder_1/operator_A_7/U2  ( .A(n2983), .B(1'b0), .Z(\adder_1/P0[7] )
         );
  AND2_X1 \adder_1/operator_A_8/U1  ( .A1(n2983), .A2(1'b0), .ZN(
        \adder_1/G0[8] ) );
  XOR2_X1 \adder_1/operator_A_8/U2  ( .A(n2983), .B(1'b0), .Z(\adder_1/P0[8] )
         );
  AND2_X1 \adder_1/operator_A_9/U1  ( .A1(n2983), .A2(1'b0), .ZN(
        \adder_1/G0[9] ) );
  XOR2_X1 \adder_1/operator_A_9/U2  ( .A(n2983), .B(1'b0), .Z(\adder_1/P0[9] )
         );
  AND2_X1 \adder_1/operator_A_10/U1  ( .A1(n2983), .A2(1'b0), .ZN(
        \adder_1/G0[10] ) );
  XOR2_X1 \adder_1/operator_A_10/U2  ( .A(n2983), .B(1'b0), .Z(
        \adder_1/P0[10] ) );
  AND2_X1 \adder_1/operator_A_11/U1  ( .A1(n2983), .A2(1'b0), .ZN(
        \adder_1/G0[11] ) );
  XOR2_X1 \adder_1/operator_A_11/U2  ( .A(n2983), .B(1'b0), .Z(
        \adder_1/P0[11] ) );
  AND2_X1 \adder_1/operator_A_12/U1  ( .A1(n2983), .A2(1'b0), .ZN(
        \adder_1/G0[12] ) );
  XOR2_X1 \adder_1/operator_A_12/U2  ( .A(n2983), .B(1'b0), .Z(
        \adder_1/P0[12] ) );
  AND2_X1 \adder_1/operator_A_13/U1  ( .A1(n2983), .A2(1'b0), .ZN(
        \adder_1/G0[13] ) );
  XOR2_X1 \adder_1/operator_A_13/U2  ( .A(n2983), .B(1'b0), .Z(
        \adder_1/P0[13] ) );
  AND2_X1 \adder_1/operator_A_14/U1  ( .A1(n2983), .A2(1'b0), .ZN(
        \adder_1/G0[14] ) );
  XOR2_X1 \adder_1/operator_A_14/U2  ( .A(n2983), .B(1'b0), .Z(
        \adder_1/P0[14] ) );
  AND2_X1 \adder_1/operator_A_15/U1  ( .A1(n2983), .A2(1'b0), .ZN(
        \adder_1/G0[15] ) );
  XOR2_X1 \adder_1/operator_A_15/U2  ( .A(n2983), .B(1'b0), .Z(
        \adder_1/P0[15] ) );
  AND2_X1 \adder_1/operator_A_16/U1  ( .A1(n2983), .A2(1'b0), .ZN(
        \adder_1/G0[16] ) );
  XOR2_X1 \adder_1/operator_A_16/U2  ( .A(n2983), .B(1'b0), .Z(
        \adder_1/P0[16] ) );
  AND2_X1 \adder_1/operator_A_17/U1  ( .A1(n2983), .A2(1'b0), .ZN(
        \adder_1/G0[17] ) );
  XOR2_X1 \adder_1/operator_A_17/U2  ( .A(n2983), .B(1'b0), .Z(
        \adder_1/P0[17] ) );
  AND2_X1 \adder_1/operator_A_18/U1  ( .A1(n2983), .A2(1'b0), .ZN(
        \adder_1/G0[18] ) );
  XOR2_X1 \adder_1/operator_A_18/U2  ( .A(n2983), .B(1'b0), .Z(
        \adder_1/P0[18] ) );
  AND2_X1 \adder_1/operator_A_19/U1  ( .A1(n3104), .A2(1'b0), .ZN(
        \adder_1/G0[19] ) );
  XOR2_X1 \adder_1/operator_A_19/U2  ( .A(n3104), .B(1'b0), .Z(
        \adder_1/P0[19] ) );
  AND2_X1 \adder_1/operator_A_20/U1  ( .A1(n3104), .A2(1'b0), .ZN(
        \adder_1/G0[20] ) );
  XOR2_X1 \adder_1/operator_A_20/U2  ( .A(n3104), .B(1'b0), .Z(
        \adder_1/P0[20] ) );
  AND2_X1 \adder_1/operator_A_21/U1  ( .A1(n3104), .A2(1'b0), .ZN(
        \adder_1/G0[21] ) );
  XOR2_X1 \adder_1/operator_A_21/U2  ( .A(n3104), .B(1'b0), .Z(
        \adder_1/P0[21] ) );
  AND2_X1 \adder_1/operator_A_22/U1  ( .A1(n3104), .A2(1'b0), .ZN(
        \adder_1/G0[22] ) );
  XOR2_X1 \adder_1/operator_A_22/U2  ( .A(n3104), .B(1'b0), .Z(
        \adder_1/P0[22] ) );
  AND2_X1 \adder_1/operator_A_23/U1  ( .A1(n3104), .A2(1'b0), .ZN(
        \adder_1/G0[23] ) );
  XOR2_X1 \adder_1/operator_A_23/U2  ( .A(n3104), .B(1'b0), .Z(
        \adder_1/P0[23] ) );
  AND2_X1 \adder_1/operator_A_24/U1  ( .A1(n2983), .A2(1'b0), .ZN(
        \adder_1/G0[24] ) );
  XOR2_X1 \adder_1/operator_A_24/U2  ( .A(n2983), .B(1'b0), .Z(
        \adder_1/P0[24] ) );
  AND2_X1 \adder_1/operator_A_25/U1  ( .A1(n2983), .A2(1'b0), .ZN(
        \adder_1/G0[25] ) );
  XOR2_X1 \adder_1/operator_A_25/U2  ( .A(n2983), .B(1'b0), .Z(
        \adder_1/P0[25] ) );
  AND2_X1 \adder_1/operator_A_26/U1  ( .A1(n2983), .A2(1'b0), .ZN(
        \adder_1/G0[26] ) );
  XOR2_X1 \adder_1/operator_A_26/U2  ( .A(n2983), .B(1'b0), .Z(
        \adder_1/P0[26] ) );
  AND2_X1 \adder_1/operator_A_27/U1  ( .A1(n2983), .A2(1'b0), .ZN(
        \adder_1/G0[27] ) );
  XOR2_X1 \adder_1/operator_A_27/U2  ( .A(n2983), .B(1'b0), .Z(
        \adder_1/P0[27] ) );
  AND2_X1 \adder_1/operator_A_28/U1  ( .A1(n2983), .A2(1'b0), .ZN(
        \adder_1/G0[28] ) );
  XOR2_X1 \adder_1/operator_A_28/U2  ( .A(n2983), .B(1'b0), .Z(
        \adder_1/P0[28] ) );
  AND2_X1 \adder_1/operator_A_29/U1  ( .A1(n2983), .A2(1'b0), .ZN(
        \adder_1/G0[29] ) );
  XOR2_X1 \adder_1/operator_A_29/U2  ( .A(n2983), .B(1'b0), .Z(
        \adder_1/P0[29] ) );
  AND2_X1 \adder_1/operator_A_30/U1  ( .A1(n2983), .A2(1'b0), .ZN(
        \adder_1/G0[30] ) );
  XOR2_X1 \adder_1/operator_A_30/U2  ( .A(n2983), .B(1'b0), .Z(
        \adder_1/P0[30] ) );
  AND2_X1 \adder_1/operator_A_31/U1  ( .A1(n2983), .A2(1'b0), .ZN(
        \adder_1/G0[31] ) );
  XOR2_X1 \adder_1/operator_A_31/U2  ( .A(n2983), .B(1'b0), .Z(
        \adder_1/P0[31] ) );
  AOI21_X1 \adder_1/operator_C_stage_1_0/U2  ( .B1(\adder_1/P0[0] ), .B2(n2983), .A(\adder_1/G0[0] ), .ZN(\adder_1/operator_C_stage_1_0/n3 ) );
  INV_X1 \adder_1/operator_C_stage_1_0/U1  ( .A(
        \adder_1/operator_C_stage_1_0/n3 ), .ZN(\adder_1/G1[0] ) );
  AOI21_X1 \adder_1/operator_B_stage_1_1/U3  ( .B1(\adder_1/G0[1] ), .B2(
        \adder_1/P0[2] ), .A(\adder_1/G0[2] ), .ZN(
        \adder_1/operator_B_stage_1_1/n3 ) );
  INV_X1 \adder_1/operator_B_stage_1_1/U2  ( .A(
        \adder_1/operator_B_stage_1_1/n3 ), .ZN(\adder_1/G1[1] ) );
  AND2_X1 \adder_1/operator_B_stage_1_1/U1  ( .A1(\adder_1/P0[1] ), .A2(
        \adder_1/P0[2] ), .ZN(\adder_1/P1[1] ) );
  AOI21_X1 \adder_1/operator_B_stage_1_2/U3  ( .B1(\adder_1/G0[3] ), .B2(
        \adder_1/P0[4] ), .A(\adder_1/G0[4] ), .ZN(
        \adder_1/operator_B_stage_1_2/n3 ) );
  INV_X1 \adder_1/operator_B_stage_1_2/U2  ( .A(
        \adder_1/operator_B_stage_1_2/n3 ), .ZN(\adder_1/G1[2] ) );
  AND2_X1 \adder_1/operator_B_stage_1_2/U1  ( .A1(\adder_1/P0[3] ), .A2(
        \adder_1/P0[4] ), .ZN(\adder_1/P1[2] ) );
  AOI21_X1 \adder_1/operator_B_stage_1_3/U3  ( .B1(\adder_1/G0[5] ), .B2(
        \adder_1/P0[6] ), .A(\adder_1/G0[6] ), .ZN(
        \adder_1/operator_B_stage_1_3/n3 ) );
  INV_X1 \adder_1/operator_B_stage_1_3/U2  ( .A(
        \adder_1/operator_B_stage_1_3/n3 ), .ZN(\adder_1/G1[3] ) );
  AND2_X1 \adder_1/operator_B_stage_1_3/U1  ( .A1(\adder_1/P0[5] ), .A2(
        \adder_1/P0[6] ), .ZN(\adder_1/P1[3] ) );
  AOI21_X1 \adder_1/operator_B_stage_1_4/U3  ( .B1(\adder_1/G0[7] ), .B2(
        \adder_1/P0[8] ), .A(\adder_1/G0[8] ), .ZN(
        \adder_1/operator_B_stage_1_4/n3 ) );
  INV_X1 \adder_1/operator_B_stage_1_4/U2  ( .A(
        \adder_1/operator_B_stage_1_4/n3 ), .ZN(\adder_1/G1[4] ) );
  AND2_X1 \adder_1/operator_B_stage_1_4/U1  ( .A1(\adder_1/P0[7] ), .A2(
        \adder_1/P0[8] ), .ZN(\adder_1/P1[4] ) );
  AOI21_X1 \adder_1/operator_B_stage_1_5/U3  ( .B1(\adder_1/G0[9] ), .B2(
        \adder_1/P0[10] ), .A(\adder_1/G0[10] ), .ZN(
        \adder_1/operator_B_stage_1_5/n3 ) );
  INV_X1 \adder_1/operator_B_stage_1_5/U2  ( .A(
        \adder_1/operator_B_stage_1_5/n3 ), .ZN(\adder_1/G1[5] ) );
  AND2_X1 \adder_1/operator_B_stage_1_5/U1  ( .A1(\adder_1/P0[9] ), .A2(
        \adder_1/P0[10] ), .ZN(\adder_1/P1[5] ) );
  AOI21_X1 \adder_1/operator_B_stage_1_6/U3  ( .B1(\adder_1/G0[11] ), .B2(
        \adder_1/P0[12] ), .A(\adder_1/G0[12] ), .ZN(
        \adder_1/operator_B_stage_1_6/n3 ) );
  INV_X1 \adder_1/operator_B_stage_1_6/U2  ( .A(
        \adder_1/operator_B_stage_1_6/n3 ), .ZN(\adder_1/G1[6] ) );
  AND2_X1 \adder_1/operator_B_stage_1_6/U1  ( .A1(\adder_1/P0[11] ), .A2(
        \adder_1/P0[12] ), .ZN(\adder_1/P1[6] ) );
  AOI21_X1 \adder_1/operator_B_stage_1_7/U3  ( .B1(\adder_1/G0[13] ), .B2(
        \adder_1/P0[14] ), .A(\adder_1/G0[14] ), .ZN(
        \adder_1/operator_B_stage_1_7/n3 ) );
  INV_X1 \adder_1/operator_B_stage_1_7/U2  ( .A(
        \adder_1/operator_B_stage_1_7/n3 ), .ZN(\adder_1/G1[7] ) );
  AND2_X1 \adder_1/operator_B_stage_1_7/U1  ( .A1(\adder_1/P0[13] ), .A2(
        \adder_1/P0[14] ), .ZN(\adder_1/P1[7] ) );
  AOI21_X1 \adder_1/operator_B_stage_1_8/U3  ( .B1(\adder_1/G0[15] ), .B2(
        \adder_1/P0[16] ), .A(\adder_1/G0[16] ), .ZN(
        \adder_1/operator_B_stage_1_8/n3 ) );
  INV_X1 \adder_1/operator_B_stage_1_8/U2  ( .A(
        \adder_1/operator_B_stage_1_8/n3 ), .ZN(\adder_1/G1[8] ) );
  AND2_X1 \adder_1/operator_B_stage_1_8/U1  ( .A1(\adder_1/P0[15] ), .A2(
        \adder_1/P0[16] ), .ZN(\adder_1/P1[8] ) );
  AOI21_X1 \adder_1/operator_B_stage_1_9/U3  ( .B1(\adder_1/G0[17] ), .B2(
        \adder_1/P0[18] ), .A(\adder_1/G0[18] ), .ZN(
        \adder_1/operator_B_stage_1_9/n3 ) );
  INV_X1 \adder_1/operator_B_stage_1_9/U2  ( .A(
        \adder_1/operator_B_stage_1_9/n3 ), .ZN(\adder_1/G1[9] ) );
  AND2_X1 \adder_1/operator_B_stage_1_9/U1  ( .A1(\adder_1/P0[17] ), .A2(
        \adder_1/P0[18] ), .ZN(\adder_1/P1[9] ) );
  AOI21_X1 \adder_1/operator_B_stage_1_10/U3  ( .B1(\adder_1/G0[19] ), .B2(
        \adder_1/P0[20] ), .A(\adder_1/G0[20] ), .ZN(
        \adder_1/operator_B_stage_1_10/n3 ) );
  INV_X1 \adder_1/operator_B_stage_1_10/U2  ( .A(
        \adder_1/operator_B_stage_1_10/n3 ), .ZN(\adder_1/G1[10] ) );
  AND2_X1 \adder_1/operator_B_stage_1_10/U1  ( .A1(\adder_1/P0[19] ), .A2(
        \adder_1/P0[20] ), .ZN(\adder_1/P1[10] ) );
  AOI21_X1 \adder_1/operator_B_stage_1_11/U3  ( .B1(\adder_1/G0[21] ), .B2(
        \adder_1/P0[22] ), .A(\adder_1/G0[22] ), .ZN(
        \adder_1/operator_B_stage_1_11/n3 ) );
  INV_X1 \adder_1/operator_B_stage_1_11/U2  ( .A(
        \adder_1/operator_B_stage_1_11/n3 ), .ZN(\adder_1/G1[11] ) );
  AND2_X1 \adder_1/operator_B_stage_1_11/U1  ( .A1(\adder_1/P0[21] ), .A2(
        \adder_1/P0[22] ), .ZN(\adder_1/P1[11] ) );
  AOI21_X1 \adder_1/operator_B_stage_1_12/U3  ( .B1(\adder_1/G0[23] ), .B2(
        \adder_1/P0[24] ), .A(\adder_1/G0[24] ), .ZN(
        \adder_1/operator_B_stage_1_12/n3 ) );
  INV_X1 \adder_1/operator_B_stage_1_12/U2  ( .A(
        \adder_1/operator_B_stage_1_12/n3 ), .ZN(\adder_1/G1[12] ) );
  AND2_X1 \adder_1/operator_B_stage_1_12/U1  ( .A1(\adder_1/P0[23] ), .A2(
        \adder_1/P0[24] ), .ZN(\adder_1/P1[12] ) );
  AOI21_X1 \adder_1/operator_B_stage_1_13/U3  ( .B1(\adder_1/G0[25] ), .B2(
        \adder_1/P0[26] ), .A(\adder_1/G0[26] ), .ZN(
        \adder_1/operator_B_stage_1_13/n3 ) );
  INV_X1 \adder_1/operator_B_stage_1_13/U2  ( .A(
        \adder_1/operator_B_stage_1_13/n3 ), .ZN(\adder_1/G1[13] ) );
  AND2_X1 \adder_1/operator_B_stage_1_13/U1  ( .A1(\adder_1/P0[25] ), .A2(
        \adder_1/P0[26] ), .ZN(\adder_1/P1[13] ) );
  AOI21_X1 \adder_1/operator_B_stage_1_14/U3  ( .B1(\adder_1/G0[27] ), .B2(
        \adder_1/P0[28] ), .A(\adder_1/G0[28] ), .ZN(
        \adder_1/operator_B_stage_1_14/n3 ) );
  INV_X1 \adder_1/operator_B_stage_1_14/U2  ( .A(
        \adder_1/operator_B_stage_1_14/n3 ), .ZN(\adder_1/G1[14] ) );
  AND2_X1 \adder_1/operator_B_stage_1_14/U1  ( .A1(\adder_1/P0[27] ), .A2(
        \adder_1/P0[28] ), .ZN(\adder_1/P1[14] ) );
  AOI21_X1 \adder_1/operator_B_stage_1_15/U3  ( .B1(\adder_1/G0[29] ), .B2(
        \adder_1/P0[30] ), .A(\adder_1/G0[30] ), .ZN(
        \adder_1/operator_B_stage_1_15/n3 ) );
  INV_X1 \adder_1/operator_B_stage_1_15/U2  ( .A(
        \adder_1/operator_B_stage_1_15/n3 ), .ZN(\adder_1/G1[15] ) );
  AND2_X1 \adder_1/operator_B_stage_1_15/U1  ( .A1(\adder_1/P0[29] ), .A2(
        \adder_1/P0[30] ), .ZN(\adder_1/P1[15] ) );
  AOI21_X1 \adder_1/operator_C_stage_2_1/U2  ( .B1(\adder_1/P1[1] ), .B2(
        \adder_1/G1[0] ), .A(\adder_1/G1[1] ), .ZN(
        \adder_1/operator_C_stage_2_1/n3 ) );
  INV_X1 \adder_1/operator_C_stage_2_1/U1  ( .A(
        \adder_1/operator_C_stage_2_1/n3 ), .ZN(\adder_1/G2[1] ) );
  AOI21_X1 \adder_1/operator_B_stage_2_2/U3  ( .B1(\adder_1/G1[1] ), .B2(
        \adder_1/P1[2] ), .A(\adder_1/G1[2] ), .ZN(
        \adder_1/operator_B_stage_2_2/n3 ) );
  INV_X1 \adder_1/operator_B_stage_2_2/U2  ( .A(
        \adder_1/operator_B_stage_2_2/n3 ), .ZN(\adder_1/G2[2] ) );
  AND2_X1 \adder_1/operator_B_stage_2_2/U1  ( .A1(\adder_1/P1[1] ), .A2(
        \adder_1/P1[2] ), .ZN(\adder_1/P2[2] ) );
  AOI21_X1 \adder_1/operator_B_stage_2_3/U3  ( .B1(\adder_1/G1[2] ), .B2(
        \adder_1/P1[3] ), .A(\adder_1/G1[3] ), .ZN(
        \adder_1/operator_B_stage_2_3/n3 ) );
  INV_X1 \adder_1/operator_B_stage_2_3/U2  ( .A(
        \adder_1/operator_B_stage_2_3/n3 ), .ZN(\adder_1/G2[3] ) );
  AND2_X1 \adder_1/operator_B_stage_2_3/U1  ( .A1(\adder_1/P1[2] ), .A2(
        \adder_1/P1[3] ), .ZN(\adder_1/P2[3] ) );
  AOI21_X1 \adder_1/operator_B_stage_2_4/U3  ( .B1(\adder_1/G1[3] ), .B2(
        \adder_1/P1[4] ), .A(\adder_1/G1[4] ), .ZN(
        \adder_1/operator_B_stage_2_4/n3 ) );
  INV_X1 \adder_1/operator_B_stage_2_4/U2  ( .A(
        \adder_1/operator_B_stage_2_4/n3 ), .ZN(\adder_1/G2[4] ) );
  AND2_X1 \adder_1/operator_B_stage_2_4/U1  ( .A1(\adder_1/P1[3] ), .A2(
        \adder_1/P1[4] ), .ZN(\adder_1/P2[4] ) );
  AOI21_X1 \adder_1/operator_B_stage_2_5/U3  ( .B1(\adder_1/G1[4] ), .B2(
        \adder_1/P1[5] ), .A(\adder_1/G1[5] ), .ZN(
        \adder_1/operator_B_stage_2_5/n3 ) );
  INV_X1 \adder_1/operator_B_stage_2_5/U2  ( .A(
        \adder_1/operator_B_stage_2_5/n3 ), .ZN(\adder_1/G2[5] ) );
  AND2_X1 \adder_1/operator_B_stage_2_5/U1  ( .A1(\adder_1/P1[4] ), .A2(
        \adder_1/P1[5] ), .ZN(\adder_1/P2[5] ) );
  AOI21_X1 \adder_1/operator_B_stage_2_6/U3  ( .B1(\adder_1/G1[5] ), .B2(
        \adder_1/P1[6] ), .A(\adder_1/G1[6] ), .ZN(
        \adder_1/operator_B_stage_2_6/n3 ) );
  INV_X1 \adder_1/operator_B_stage_2_6/U2  ( .A(
        \adder_1/operator_B_stage_2_6/n3 ), .ZN(\adder_1/G2[6] ) );
  AND2_X1 \adder_1/operator_B_stage_2_6/U1  ( .A1(\adder_1/P1[5] ), .A2(
        \adder_1/P1[6] ), .ZN(\adder_1/P2[6] ) );
  AOI21_X1 \adder_1/operator_B_stage_2_7/U3  ( .B1(\adder_1/G1[6] ), .B2(
        \adder_1/P1[7] ), .A(\adder_1/G1[7] ), .ZN(
        \adder_1/operator_B_stage_2_7/n3 ) );
  INV_X1 \adder_1/operator_B_stage_2_7/U2  ( .A(
        \adder_1/operator_B_stage_2_7/n3 ), .ZN(\adder_1/G2[7] ) );
  AND2_X1 \adder_1/operator_B_stage_2_7/U1  ( .A1(\adder_1/P1[6] ), .A2(
        \adder_1/P1[7] ), .ZN(\adder_1/P2[7] ) );
  AOI21_X1 \adder_1/operator_B_stage_2_8/U3  ( .B1(\adder_1/G1[7] ), .B2(
        \adder_1/P1[8] ), .A(\adder_1/G1[8] ), .ZN(
        \adder_1/operator_B_stage_2_8/n3 ) );
  INV_X1 \adder_1/operator_B_stage_2_8/U2  ( .A(
        \adder_1/operator_B_stage_2_8/n3 ), .ZN(\adder_1/G2[8] ) );
  AND2_X1 \adder_1/operator_B_stage_2_8/U1  ( .A1(\adder_1/P1[7] ), .A2(
        \adder_1/P1[8] ), .ZN(\adder_1/P2[8] ) );
  AOI21_X1 \adder_1/operator_B_stage_2_9/U3  ( .B1(\adder_1/G1[8] ), .B2(
        \adder_1/P1[9] ), .A(\adder_1/G1[9] ), .ZN(
        \adder_1/operator_B_stage_2_9/n3 ) );
  INV_X1 \adder_1/operator_B_stage_2_9/U2  ( .A(
        \adder_1/operator_B_stage_2_9/n3 ), .ZN(\adder_1/G2[9] ) );
  AND2_X1 \adder_1/operator_B_stage_2_9/U1  ( .A1(\adder_1/P1[8] ), .A2(
        \adder_1/P1[9] ), .ZN(\adder_1/P2[9] ) );
  AOI21_X1 \adder_1/operator_B_stage_2_10/U3  ( .B1(\adder_1/G1[9] ), .B2(
        \adder_1/P1[10] ), .A(\adder_1/G1[10] ), .ZN(
        \adder_1/operator_B_stage_2_10/n3 ) );
  INV_X1 \adder_1/operator_B_stage_2_10/U2  ( .A(
        \adder_1/operator_B_stage_2_10/n3 ), .ZN(\adder_1/G2[10] ) );
  AND2_X1 \adder_1/operator_B_stage_2_10/U1  ( .A1(\adder_1/P1[9] ), .A2(
        \adder_1/P1[10] ), .ZN(\adder_1/P2[10] ) );
  AOI21_X1 \adder_1/operator_B_stage_2_11/U3  ( .B1(\adder_1/G1[10] ), .B2(
        \adder_1/P1[11] ), .A(\adder_1/G1[11] ), .ZN(
        \adder_1/operator_B_stage_2_11/n3 ) );
  INV_X1 \adder_1/operator_B_stage_2_11/U2  ( .A(
        \adder_1/operator_B_stage_2_11/n3 ), .ZN(\adder_1/G2[11] ) );
  AND2_X1 \adder_1/operator_B_stage_2_11/U1  ( .A1(\adder_1/P1[10] ), .A2(
        \adder_1/P1[11] ), .ZN(\adder_1/P2[11] ) );
  AOI21_X1 \adder_1/operator_B_stage_2_12/U3  ( .B1(\adder_1/G1[11] ), .B2(
        \adder_1/P1[12] ), .A(\adder_1/G1[12] ), .ZN(
        \adder_1/operator_B_stage_2_12/n3 ) );
  INV_X1 \adder_1/operator_B_stage_2_12/U2  ( .A(
        \adder_1/operator_B_stage_2_12/n3 ), .ZN(\adder_1/G2[12] ) );
  AND2_X1 \adder_1/operator_B_stage_2_12/U1  ( .A1(\adder_1/P1[11] ), .A2(
        \adder_1/P1[12] ), .ZN(\adder_1/P2[12] ) );
  AOI21_X1 \adder_1/operator_B_stage_2_13/U3  ( .B1(\adder_1/G1[12] ), .B2(
        \adder_1/P1[13] ), .A(\adder_1/G1[13] ), .ZN(
        \adder_1/operator_B_stage_2_13/n3 ) );
  INV_X1 \adder_1/operator_B_stage_2_13/U2  ( .A(
        \adder_1/operator_B_stage_2_13/n3 ), .ZN(\adder_1/G2[13] ) );
  AND2_X1 \adder_1/operator_B_stage_2_13/U1  ( .A1(\adder_1/P1[12] ), .A2(
        \adder_1/P1[13] ), .ZN(\adder_1/P2[13] ) );
  AOI21_X1 \adder_1/operator_B_stage_2_14/U3  ( .B1(\adder_1/G1[13] ), .B2(
        \adder_1/P1[14] ), .A(\adder_1/G1[14] ), .ZN(
        \adder_1/operator_B_stage_2_14/n3 ) );
  AND2_X1 \adder_1/operator_B_stage_2_14/U2  ( .A1(\adder_1/P1[13] ), .A2(
        \adder_1/P1[14] ), .ZN(\adder_1/P2[14] ) );
  INV_X1 \adder_1/operator_B_stage_2_14/U1  ( .A(
        \adder_1/operator_B_stage_2_14/n3 ), .ZN(\adder_1/G2[14] ) );
  AOI21_X1 \adder_1/operator_B_stage_2_15/U3  ( .B1(\adder_1/G1[14] ), .B2(
        \adder_1/P1[15] ), .A(\adder_1/G1[15] ), .ZN(
        \adder_1/operator_B_stage_2_15/n3 ) );
  INV_X1 \adder_1/operator_B_stage_2_15/U2  ( .A(
        \adder_1/operator_B_stage_2_15/n3 ), .ZN(\adder_1/G2[15] ) );
  AND2_X1 \adder_1/operator_B_stage_2_15/U1  ( .A1(\adder_1/P1[14] ), .A2(
        \adder_1/P1[15] ), .ZN(\adder_1/P2[15] ) );
  AOI21_X1 \adder_1/operator_C_stage_3_2/U2  ( .B1(\adder_1/P2[2] ), .B2(
        \adder_1/G1[0] ), .A(\adder_1/G2[2] ), .ZN(
        \adder_1/operator_C_stage_3_2/n3 ) );
  INV_X1 \adder_1/operator_C_stage_3_2/U1  ( .A(
        \adder_1/operator_C_stage_3_2/n3 ), .ZN(\adder_1/G3[2] ) );
  AOI21_X1 \adder_1/operator_C_stage_3_3/U2  ( .B1(\adder_1/P2[3] ), .B2(
        \adder_1/G2[1] ), .A(\adder_1/G2[3] ), .ZN(
        \adder_1/operator_C_stage_3_3/n3 ) );
  INV_X1 \adder_1/operator_C_stage_3_3/U1  ( .A(
        \adder_1/operator_C_stage_3_3/n3 ), .ZN(\adder_1/G3[3] ) );
  AOI21_X1 \adder_1/operator_B_stage_3_4/U3  ( .B1(\adder_1/G2[2] ), .B2(
        \adder_1/P2[4] ), .A(\adder_1/G2[4] ), .ZN(
        \adder_1/operator_B_stage_3_4/n3 ) );
  INV_X1 \adder_1/operator_B_stage_3_4/U2  ( .A(
        \adder_1/operator_B_stage_3_4/n3 ), .ZN(\adder_1/G3[4] ) );
  AND2_X1 \adder_1/operator_B_stage_3_4/U1  ( .A1(\adder_1/P2[2] ), .A2(
        \adder_1/P2[4] ), .ZN(\adder_1/P3[4] ) );
  AOI21_X1 \adder_1/operator_B_stage_3_5/U3  ( .B1(\adder_1/G2[3] ), .B2(
        \adder_1/P2[5] ), .A(\adder_1/G2[5] ), .ZN(
        \adder_1/operator_B_stage_3_5/n3 ) );
  INV_X1 \adder_1/operator_B_stage_3_5/U2  ( .A(
        \adder_1/operator_B_stage_3_5/n3 ), .ZN(\adder_1/G3[5] ) );
  AND2_X1 \adder_1/operator_B_stage_3_5/U1  ( .A1(\adder_1/P2[3] ), .A2(
        \adder_1/P2[5] ), .ZN(\adder_1/P3[5] ) );
  AOI21_X1 \adder_1/operator_B_stage_3_6/U3  ( .B1(\adder_1/G2[4] ), .B2(
        \adder_1/P2[6] ), .A(\adder_1/G2[6] ), .ZN(
        \adder_1/operator_B_stage_3_6/n3 ) );
  INV_X1 \adder_1/operator_B_stage_3_6/U2  ( .A(
        \adder_1/operator_B_stage_3_6/n3 ), .ZN(\adder_1/G3[6] ) );
  AND2_X1 \adder_1/operator_B_stage_3_6/U1  ( .A1(\adder_1/P2[4] ), .A2(
        \adder_1/P2[6] ), .ZN(\adder_1/P3[6] ) );
  AOI21_X1 \adder_1/operator_B_stage_3_7/U3  ( .B1(\adder_1/G2[5] ), .B2(
        \adder_1/P2[7] ), .A(\adder_1/G2[7] ), .ZN(
        \adder_1/operator_B_stage_3_7/n3 ) );
  INV_X1 \adder_1/operator_B_stage_3_7/U2  ( .A(
        \adder_1/operator_B_stage_3_7/n3 ), .ZN(\adder_1/G3[7] ) );
  AND2_X1 \adder_1/operator_B_stage_3_7/U1  ( .A1(\adder_1/P2[5] ), .A2(
        \adder_1/P2[7] ), .ZN(\adder_1/P3[7] ) );
  AOI21_X1 \adder_1/operator_B_stage_3_8/U3  ( .B1(\adder_1/G2[6] ), .B2(
        \adder_1/P2[8] ), .A(\adder_1/G2[8] ), .ZN(
        \adder_1/operator_B_stage_3_8/n3 ) );
  INV_X1 \adder_1/operator_B_stage_3_8/U2  ( .A(
        \adder_1/operator_B_stage_3_8/n3 ), .ZN(\adder_1/G3[8] ) );
  AND2_X1 \adder_1/operator_B_stage_3_8/U1  ( .A1(\adder_1/P2[6] ), .A2(
        \adder_1/P2[8] ), .ZN(\adder_1/P3[8] ) );
  AOI21_X1 \adder_1/operator_B_stage_3_9/U3  ( .B1(\adder_1/G2[7] ), .B2(
        \adder_1/P2[9] ), .A(\adder_1/G2[9] ), .ZN(
        \adder_1/operator_B_stage_3_9/n3 ) );
  INV_X1 \adder_1/operator_B_stage_3_9/U2  ( .A(
        \adder_1/operator_B_stage_3_9/n3 ), .ZN(\adder_1/G3[9] ) );
  AND2_X1 \adder_1/operator_B_stage_3_9/U1  ( .A1(\adder_1/P2[7] ), .A2(
        \adder_1/P2[9] ), .ZN(\adder_1/P3[9] ) );
  AOI21_X1 \adder_1/operator_B_stage_3_10/U3  ( .B1(\adder_1/G2[8] ), .B2(
        \adder_1/P2[10] ), .A(\adder_1/G2[10] ), .ZN(
        \adder_1/operator_B_stage_3_10/n3 ) );
  INV_X1 \adder_1/operator_B_stage_3_10/U2  ( .A(
        \adder_1/operator_B_stage_3_10/n3 ), .ZN(\adder_1/G3[10] ) );
  AND2_X1 \adder_1/operator_B_stage_3_10/U1  ( .A1(\adder_1/P2[8] ), .A2(
        \adder_1/P2[10] ), .ZN(\adder_1/P3[10] ) );
  AOI21_X1 \adder_1/operator_B_stage_3_11/U3  ( .B1(\adder_1/G2[9] ), .B2(
        \adder_1/P2[11] ), .A(\adder_1/G2[11] ), .ZN(
        \adder_1/operator_B_stage_3_11/n3 ) );
  INV_X1 \adder_1/operator_B_stage_3_11/U2  ( .A(
        \adder_1/operator_B_stage_3_11/n3 ), .ZN(\adder_1/G3[11] ) );
  AND2_X1 \adder_1/operator_B_stage_3_11/U1  ( .A1(\adder_1/P2[9] ), .A2(
        \adder_1/P2[11] ), .ZN(\adder_1/P3[11] ) );
  AOI21_X1 \adder_1/operator_B_stage_3_12/U3  ( .B1(\adder_1/G2[10] ), .B2(
        \adder_1/P2[12] ), .A(\adder_1/G2[12] ), .ZN(
        \adder_1/operator_B_stage_3_12/n3 ) );
  INV_X1 \adder_1/operator_B_stage_3_12/U2  ( .A(
        \adder_1/operator_B_stage_3_12/n3 ), .ZN(\adder_1/G3[12] ) );
  AND2_X1 \adder_1/operator_B_stage_3_12/U1  ( .A1(\adder_1/P2[10] ), .A2(
        \adder_1/P2[12] ), .ZN(\adder_1/P3[12] ) );
  AOI21_X1 \adder_1/operator_B_stage_3_13/U3  ( .B1(\adder_1/G2[11] ), .B2(
        \adder_1/P2[13] ), .A(\adder_1/G2[13] ), .ZN(
        \adder_1/operator_B_stage_3_13/n3 ) );
  INV_X1 \adder_1/operator_B_stage_3_13/U2  ( .A(
        \adder_1/operator_B_stage_3_13/n3 ), .ZN(\adder_1/G3[13] ) );
  AND2_X1 \adder_1/operator_B_stage_3_13/U1  ( .A1(\adder_1/P2[11] ), .A2(
        \adder_1/P2[13] ), .ZN(\adder_1/P3[13] ) );
  AOI21_X1 \adder_1/operator_B_stage_3_14/U3  ( .B1(\adder_1/G2[12] ), .B2(
        \adder_1/P2[14] ), .A(\adder_1/G2[14] ), .ZN(
        \adder_1/operator_B_stage_3_14/n3 ) );
  INV_X1 \adder_1/operator_B_stage_3_14/U2  ( .A(
        \adder_1/operator_B_stage_3_14/n3 ), .ZN(\adder_1/G3[14] ) );
  AND2_X1 \adder_1/operator_B_stage_3_14/U1  ( .A1(\adder_1/P2[12] ), .A2(
        \adder_1/P2[14] ), .ZN(\adder_1/P3[14] ) );
  AOI21_X1 \adder_1/operator_B_stage_3_15/U3  ( .B1(\adder_1/G2[13] ), .B2(
        \adder_1/P2[15] ), .A(\adder_1/G2[15] ), .ZN(
        \adder_1/operator_B_stage_3_15/n3 ) );
  INV_X1 \adder_1/operator_B_stage_3_15/U2  ( .A(
        \adder_1/operator_B_stage_3_15/n3 ), .ZN(\adder_1/G3[15] ) );
  AND2_X1 \adder_1/operator_B_stage_3_15/U1  ( .A1(\adder_1/P2[13] ), .A2(
        \adder_1/P2[15] ), .ZN(\adder_1/P3[15] ) );
  AOI21_X1 \adder_1/operator_C_stage_4_4/U2  ( .B1(\adder_1/P3[4] ), .B2(
        \adder_1/G1[0] ), .A(\adder_1/G3[4] ), .ZN(
        \adder_1/operator_C_stage_4_4/n3 ) );
  INV_X1 \adder_1/operator_C_stage_4_4/U1  ( .A(
        \adder_1/operator_C_stage_4_4/n3 ), .ZN(\adder_1/G4[4] ) );
  AOI21_X1 \adder_1/operator_C_stage_4_5/U2  ( .B1(\adder_1/P3[5] ), .B2(
        \adder_1/G2[1] ), .A(\adder_1/G3[5] ), .ZN(
        \adder_1/operator_C_stage_4_5/n3 ) );
  INV_X1 \adder_1/operator_C_stage_4_5/U1  ( .A(
        \adder_1/operator_C_stage_4_5/n3 ), .ZN(\adder_1/G4[5] ) );
  AOI21_X1 \adder_1/operator_C_stage_4_6/U2  ( .B1(\adder_1/P3[6] ), .B2(
        \adder_1/G3[2] ), .A(\adder_1/G3[6] ), .ZN(
        \adder_1/operator_C_stage_4_6/n3 ) );
  INV_X1 \adder_1/operator_C_stage_4_6/U1  ( .A(
        \adder_1/operator_C_stage_4_6/n3 ), .ZN(\adder_1/G4[6] ) );
  AOI21_X1 \adder_1/operator_C_stage_4_7/U2  ( .B1(\adder_1/P3[7] ), .B2(
        \adder_1/G3[3] ), .A(\adder_1/G3[7] ), .ZN(
        \adder_1/operator_C_stage_4_7/n3 ) );
  INV_X1 \adder_1/operator_C_stage_4_7/U1  ( .A(
        \adder_1/operator_C_stage_4_7/n3 ), .ZN(\adder_1/G4[7] ) );
  AND2_X1 \adder_1/operator_B_stage_4_8/U3  ( .A1(\adder_1/P3[4] ), .A2(
        \adder_1/P3[8] ), .ZN(\adder_1/P4 [8]) );
  INV_X1 \adder_1/operator_B_stage_4_8/U2  ( .A(
        \adder_1/operator_B_stage_4_8/n3 ), .ZN(\adder_1/G4[8] ) );
  AOI21_X1 \adder_1/operator_B_stage_4_8/U1  ( .B1(\adder_1/G3[4] ), .B2(
        \adder_1/P3[8] ), .A(\adder_1/G3[8] ), .ZN(
        \adder_1/operator_B_stage_4_8/n3 ) );
  AND2_X1 \adder_1/operator_B_stage_4_9/U3  ( .A1(\adder_1/P3[5] ), .A2(
        \adder_1/P3[9] ), .ZN(\adder_1/P4 [9]) );
  INV_X1 \adder_1/operator_B_stage_4_9/U2  ( .A(
        \adder_1/operator_B_stage_4_9/n3 ), .ZN(\adder_1/G4[9] ) );
  AOI21_X1 \adder_1/operator_B_stage_4_9/U1  ( .B1(\adder_1/G3[5] ), .B2(
        \adder_1/P3[9] ), .A(\adder_1/G3[9] ), .ZN(
        \adder_1/operator_B_stage_4_9/n3 ) );
  AND2_X1 \adder_1/operator_B_stage_4_10/U3  ( .A1(\adder_1/P3[6] ), .A2(
        \adder_1/P3[10] ), .ZN(\adder_1/P4 [10]) );
  INV_X1 \adder_1/operator_B_stage_4_10/U2  ( .A(
        \adder_1/operator_B_stage_4_10/n3 ), .ZN(\adder_1/G4[10] ) );
  AOI21_X1 \adder_1/operator_B_stage_4_10/U1  ( .B1(\adder_1/G3[6] ), .B2(
        \adder_1/P3[10] ), .A(\adder_1/G3[10] ), .ZN(
        \adder_1/operator_B_stage_4_10/n3 ) );
  AND2_X1 \adder_1/operator_B_stage_4_11/U3  ( .A1(\adder_1/P3[7] ), .A2(
        \adder_1/P3[11] ), .ZN(\adder_1/P4 [11]) );
  INV_X1 \adder_1/operator_B_stage_4_11/U2  ( .A(
        \adder_1/operator_B_stage_4_11/n3 ), .ZN(\adder_1/G4[11] ) );
  AOI21_X1 \adder_1/operator_B_stage_4_11/U1  ( .B1(\adder_1/G3[7] ), .B2(
        \adder_1/P3[11] ), .A(\adder_1/G3[11] ), .ZN(
        \adder_1/operator_B_stage_4_11/n3 ) );
  AND2_X1 \adder_1/operator_B_stage_4_12/U3  ( .A1(\adder_1/P3[8] ), .A2(
        \adder_1/P3[12] ), .ZN(\adder_1/P4 [12]) );
  INV_X1 \adder_1/operator_B_stage_4_12/U2  ( .A(
        \adder_1/operator_B_stage_4_12/n3 ), .ZN(\adder_1/G4[12] ) );
  AOI21_X1 \adder_1/operator_B_stage_4_12/U1  ( .B1(\adder_1/G3[8] ), .B2(
        \adder_1/P3[12] ), .A(\adder_1/G3[12] ), .ZN(
        \adder_1/operator_B_stage_4_12/n3 ) );
  AOI21_X1 \adder_1/operator_B_stage_4_13/U3  ( .B1(\adder_1/G3[9] ), .B2(
        \adder_1/P3[13] ), .A(\adder_1/G3[13] ), .ZN(
        \adder_1/operator_B_stage_4_13/n3 ) );
  AND2_X1 \adder_1/operator_B_stage_4_13/U2  ( .A1(\adder_1/P3[9] ), .A2(
        \adder_1/P3[13] ), .ZN(\adder_1/P4 [13]) );
  INV_X1 \adder_1/operator_B_stage_4_13/U1  ( .A(
        \adder_1/operator_B_stage_4_13/n3 ), .ZN(\adder_1/G4[13] ) );
  AOI21_X1 \adder_1/operator_B_stage_4_14/U3  ( .B1(\adder_1/G3[10] ), .B2(
        \adder_1/P3[14] ), .A(\adder_1/G3[14] ), .ZN(
        \adder_1/operator_B_stage_4_14/n3 ) );
  AND2_X1 \adder_1/operator_B_stage_4_14/U2  ( .A1(\adder_1/P3[10] ), .A2(
        \adder_1/P3[14] ), .ZN(\adder_1/P4 [14]) );
  INV_X1 \adder_1/operator_B_stage_4_14/U1  ( .A(
        \adder_1/operator_B_stage_4_14/n3 ), .ZN(\adder_1/G4[14] ) );
  AOI21_X1 \adder_1/operator_B_stage_4_15/U3  ( .B1(\adder_1/G3[11] ), .B2(
        \adder_1/P3[15] ), .A(\adder_1/G3[15] ), .ZN(
        \adder_1/operator_B_stage_4_15/n3 ) );
  AND2_X1 \adder_1/operator_B_stage_4_15/U2  ( .A1(\adder_1/P3[11] ), .A2(
        \adder_1/P3[15] ), .ZN(\adder_1/P4 [15]) );
  INV_X1 \adder_1/operator_B_stage_4_15/U1  ( .A(
        \adder_1/operator_B_stage_4_15/n3 ), .ZN(\adder_1/G4[15] ) );
  AOI21_X1 \adder_1/operator_C_stage_5_8/U2  ( .B1(\adder_1/P4 [8]), .B2(
        \adder_1/G1[0] ), .A(\adder_1/G4[8] ), .ZN(
        \adder_1/operator_C_stage_5_8/n3 ) );
  INV_X1 \adder_1/operator_C_stage_5_8/U1  ( .A(
        \adder_1/operator_C_stage_5_8/n3 ), .ZN(\adder_1/G5[8] ) );
  AOI21_X1 \adder_1/operator_C_stage_5_9/U2  ( .B1(\adder_1/P4 [9]), .B2(
        \adder_1/G2[1] ), .A(\adder_1/G4[9] ), .ZN(
        \adder_1/operator_C_stage_5_9/n3 ) );
  INV_X1 \adder_1/operator_C_stage_5_9/U1  ( .A(
        \adder_1/operator_C_stage_5_9/n3 ), .ZN(\adder_1/G5[9] ) );
  AOI21_X1 \adder_1/operator_C_stage_5_10/U2  ( .B1(\adder_1/P4 [10]), .B2(
        \adder_1/G3[2] ), .A(\adder_1/G4[10] ), .ZN(
        \adder_1/operator_C_stage_5_10/n3 ) );
  INV_X1 \adder_1/operator_C_stage_5_10/U1  ( .A(
        \adder_1/operator_C_stage_5_10/n3 ), .ZN(\adder_1/G5[10] ) );
  AOI21_X1 \adder_1/operator_C_stage_5_11/U2  ( .B1(\adder_1/P4 [11]), .B2(
        \adder_1/G3[3] ), .A(\adder_1/G4[11] ), .ZN(
        \adder_1/operator_C_stage_5_11/n3 ) );
  INV_X1 \adder_1/operator_C_stage_5_11/U1  ( .A(
        \adder_1/operator_C_stage_5_11/n3 ), .ZN(\adder_1/G5[11] ) );
  AOI21_X1 \adder_1/operator_C_stage_5_12/U2  ( .B1(\adder_1/P4 [12]), .B2(
        \adder_1/G4[4] ), .A(\adder_1/G4[12] ), .ZN(
        \adder_1/operator_C_stage_5_12/n3 ) );
  INV_X1 \adder_1/operator_C_stage_5_12/U1  ( .A(
        \adder_1/operator_C_stage_5_12/n3 ), .ZN(\adder_1/G5[12] ) );
  AOI21_X1 \adder_1/operator_C_stage_5_13/U2  ( .B1(\adder_1/P4 [13]), .B2(
        \adder_1/G4[5] ), .A(\adder_1/G4[13] ), .ZN(
        \adder_1/operator_C_stage_5_13/n3 ) );
  INV_X1 \adder_1/operator_C_stage_5_13/U1  ( .A(
        \adder_1/operator_C_stage_5_13/n3 ), .ZN(\adder_1/G5[13] ) );
  AOI21_X1 \adder_1/operator_C_stage_5_14/U2  ( .B1(\adder_1/P4 [14]), .B2(
        \adder_1/G4[6] ), .A(\adder_1/G4[14] ), .ZN(
        \adder_1/operator_C_stage_5_14/n3 ) );
  INV_X1 \adder_1/operator_C_stage_5_14/U1  ( .A(
        \adder_1/operator_C_stage_5_14/n3 ), .ZN(\adder_1/G5[14] ) );
  AOI21_X1 \adder_1/operator_C_stage_5_15/U2  ( .B1(\adder_1/P4 [15]), .B2(
        \adder_1/G4[7] ), .A(\adder_1/G4[15] ), .ZN(
        \adder_1/operator_C_stage_5_15/n3 ) );
  INV_X1 \adder_1/operator_C_stage_5_15/U1  ( .A(
        \adder_1/operator_C_stage_5_15/n3 ), .ZN(\adder_1/G5[15] ) );
  INV_X1 \adder_1/operator_C_stage_6_0/U2  ( .A(
        \adder_1/operator_C_stage_6_0/n3 ), .ZN(\adder_1/G6_1 ) );
  AOI21_X1 \adder_1/operator_C_stage_6_0/U1  ( .B1(\adder_1/P0[1] ), .B2(
        \adder_1/G1[0] ), .A(\adder_1/G0[1] ), .ZN(
        \adder_1/operator_C_stage_6_0/n3 ) );
  INV_X1 \adder_1/operator_C_stage_6_1/U2  ( .A(
        \adder_1/operator_C_stage_6_1/n3 ), .ZN(\adder_1/G6_3 ) );
  AOI21_X1 \adder_1/operator_C_stage_6_1/U1  ( .B1(\adder_1/P0[3] ), .B2(
        \adder_1/G2[1] ), .A(\adder_1/G0[3] ), .ZN(
        \adder_1/operator_C_stage_6_1/n3 ) );
  AOI21_X1 \adder_1/operator_C_stage_6_2/U2  ( .B1(\adder_1/P0[5] ), .B2(
        \adder_1/G3[2] ), .A(\adder_1/G0[5] ), .ZN(
        \adder_1/operator_C_stage_6_2/n3 ) );
  INV_X1 \adder_1/operator_C_stage_6_2/U1  ( .A(
        \adder_1/operator_C_stage_6_2/n3 ), .ZN(\adder_1/G6_5 ) );
  AOI21_X1 \adder_1/operator_C_stage_6_3/U2  ( .B1(\adder_1/P0[7] ), .B2(
        \adder_1/G3[3] ), .A(\adder_1/G0[7] ), .ZN(
        \adder_1/operator_C_stage_6_3/n3 ) );
  INV_X1 \adder_1/operator_C_stage_6_3/U1  ( .A(
        \adder_1/operator_C_stage_6_3/n3 ), .ZN(\adder_1/G6_7 ) );
  AOI21_X1 \adder_1/operator_C_stage_6_4/U2  ( .B1(\adder_1/P0[9] ), .B2(
        \adder_1/G4[4] ), .A(\adder_1/G0[9] ), .ZN(
        \adder_1/operator_C_stage_6_4/n3 ) );
  INV_X1 \adder_1/operator_C_stage_6_4/U1  ( .A(
        \adder_1/operator_C_stage_6_4/n3 ), .ZN(\adder_1/G6_9 ) );
  AOI21_X1 \adder_1/operator_C_stage_6_5/U2  ( .B1(\adder_1/P0[11] ), .B2(
        \adder_1/G4[5] ), .A(\adder_1/G0[11] ), .ZN(
        \adder_1/operator_C_stage_6_5/n3 ) );
  INV_X1 \adder_1/operator_C_stage_6_5/U1  ( .A(
        \adder_1/operator_C_stage_6_5/n3 ), .ZN(\adder_1/G6_11 ) );
  AOI21_X1 \adder_1/operator_C_stage_6_6/U2  ( .B1(\adder_1/P0[13] ), .B2(
        \adder_1/G4[6] ), .A(\adder_1/G0[13] ), .ZN(
        \adder_1/operator_C_stage_6_6/n3 ) );
  INV_X1 \adder_1/operator_C_stage_6_6/U1  ( .A(
        \adder_1/operator_C_stage_6_6/n3 ), .ZN(\adder_1/G6_13 ) );
  AOI21_X1 \adder_1/operator_C_stage_6_7/U2  ( .B1(\adder_1/P0[15] ), .B2(
        \adder_1/G4[7] ), .A(\adder_1/G0[15] ), .ZN(
        \adder_1/operator_C_stage_6_7/n3 ) );
  INV_X1 \adder_1/operator_C_stage_6_7/U1  ( .A(
        \adder_1/operator_C_stage_6_7/n3 ), .ZN(\adder_1/G6_15 ) );
  AOI21_X1 \adder_1/operator_C_stage_6_8/U2  ( .B1(\adder_1/P0[17] ), .B2(
        \adder_1/G5[8] ), .A(\adder_1/G0[17] ), .ZN(
        \adder_1/operator_C_stage_6_8/n3 ) );
  INV_X1 \adder_1/operator_C_stage_6_8/U1  ( .A(
        \adder_1/operator_C_stage_6_8/n3 ), .ZN(\adder_1/G6_17 ) );
  AOI21_X1 \adder_1/operator_C_stage_6_9/U2  ( .B1(\adder_1/P0[19] ), .B2(
        \adder_1/G5[9] ), .A(\adder_1/G0[19] ), .ZN(
        \adder_1/operator_C_stage_6_9/n3 ) );
  INV_X1 \adder_1/operator_C_stage_6_9/U1  ( .A(
        \adder_1/operator_C_stage_6_9/n3 ), .ZN(\adder_1/G6_19 ) );
  AOI21_X1 \adder_1/operator_C_stage_6_10/U2  ( .B1(\adder_1/P0[21] ), .B2(
        \adder_1/G5[10] ), .A(\adder_1/G0[21] ), .ZN(
        \adder_1/operator_C_stage_6_10/n3 ) );
  INV_X1 \adder_1/operator_C_stage_6_10/U1  ( .A(
        \adder_1/operator_C_stage_6_10/n3 ), .ZN(\adder_1/G6_21 ) );
  AOI21_X1 \adder_1/operator_C_stage_6_11/U2  ( .B1(\adder_1/P0[23] ), .B2(
        \adder_1/G5[11] ), .A(\adder_1/G0[23] ), .ZN(
        \adder_1/operator_C_stage_6_11/n3 ) );
  INV_X1 \adder_1/operator_C_stage_6_11/U1  ( .A(
        \adder_1/operator_C_stage_6_11/n3 ), .ZN(\adder_1/G6_23 ) );
  AOI21_X1 \adder_1/operator_C_stage_6_12/U2  ( .B1(\adder_1/P0[25] ), .B2(
        \adder_1/G5[12] ), .A(\adder_1/G0[25] ), .ZN(
        \adder_1/operator_C_stage_6_12/n3 ) );
  INV_X1 \adder_1/operator_C_stage_6_12/U1  ( .A(
        \adder_1/operator_C_stage_6_12/n3 ), .ZN(\adder_1/G6_25 ) );
  AOI21_X1 \adder_1/operator_C_stage_6_13/U2  ( .B1(\adder_1/P0[27] ), .B2(
        \adder_1/G5[13] ), .A(\adder_1/G0[27] ), .ZN(
        \adder_1/operator_C_stage_6_13/n3 ) );
  INV_X1 \adder_1/operator_C_stage_6_13/U1  ( .A(
        \adder_1/operator_C_stage_6_13/n3 ), .ZN(\adder_1/G6_27 ) );
  AOI21_X1 \adder_1/operator_C_stage_6_14/U2  ( .B1(\adder_1/P0[29] ), .B2(
        \adder_1/G5[14] ), .A(\adder_1/G0[29] ), .ZN(
        \adder_1/operator_C_stage_6_14/n3 ) );
  INV_X1 \adder_1/operator_C_stage_6_14/U1  ( .A(
        \adder_1/operator_C_stage_6_14/n3 ), .ZN(\adder_1/G6_29_ ) );
  AOI21_X1 \adder_1/operator_C_stage_6_15/U2  ( .B1(\adder_1/P0[31] ), .B2(
        \adder_1/G5[15] ), .A(\adder_1/G0[31] ), .ZN(
        \adder_1/operator_C_stage_6_15/n3 ) );
  INV_X1 \adder_1/operator_C_stage_6_15/U1  ( .A(
        \adder_1/operator_C_stage_6_15/n3 ), .ZN(\adder_1/o_c ) );
  BUF_X1 \sra_198/U249  ( .A(PR_1[31]), .Z(N295) );
  INV_X1 \sra_198/U248  ( .A(PR_1[27]), .ZN(\sra_198/n286 ) );
  INV_X1 \sra_198/U247  ( .A(PR_1[30]), .ZN(\sra_198/n289 ) );
  INV_X1 \sra_198/U246  ( .A(PR_1[3]), .ZN(\sra_198/n262 ) );
  INV_X1 \sra_198/U245  ( .A(PR_1[4]), .ZN(\sra_198/n263 ) );
  INV_X1 \sra_198/U244  ( .A(PR_1[5]), .ZN(\sra_198/n264 ) );
  INV_X1 \sra_198/U243  ( .A(PR_1[14]), .ZN(\sra_198/n273 ) );
  INV_X1 \sra_198/U242  ( .A(PR_1[15]), .ZN(\sra_198/n274 ) );
  INV_X1 \sra_198/U241  ( .A(PR_1[11]), .ZN(\sra_198/n270 ) );
  INV_X1 \sra_198/U240  ( .A(PR_1[19]), .ZN(\sra_198/n278 ) );
  INV_X1 \sra_198/U239  ( .A(PR_1[18]), .ZN(\sra_198/n277 ) );
  INV_X1 \sra_198/U238  ( .A(PR_1[20]), .ZN(\sra_198/n279 ) );
  INV_X1 \sra_198/U237  ( .A(PR_1[16]), .ZN(\sra_198/n275 ) );
  INV_X1 \sra_198/U236  ( .A(PR_1[12]), .ZN(\sra_198/n271 ) );
  INV_X1 \sra_198/U235  ( .A(PR_1[21]), .ZN(\sra_198/n280 ) );
  INV_X1 \sra_198/U234  ( .A(PR_1[22]), .ZN(\sra_198/n281 ) );
  INV_X1 \sra_198/U233  ( .A(PR_1[23]), .ZN(\sra_198/n282 ) );
  INV_X1 \sra_198/U232  ( .A(PR_1[24]), .ZN(\sra_198/n283 ) );
  INV_X1 \sra_198/U231  ( .A(PR_1[13]), .ZN(\sra_198/n272 ) );
  INV_X1 \sra_198/U230  ( .A(PR_1[17]), .ZN(\sra_198/n276 ) );
  INV_X1 \sra_198/U229  ( .A(PR_1[25]), .ZN(\sra_198/n284 ) );
  INV_X1 \sra_198/U228  ( .A(PR_1[26]), .ZN(\sra_198/n285 ) );
  INV_X1 \sra_198/U227  ( .A(PR_1[28]), .ZN(\sra_198/n287 ) );
  INV_X1 \sra_198/U225  ( .A(PR_1[6]), .ZN(\sra_198/n265 ) );
  INV_X1 \sra_198/U224  ( .A(PR_1[7]), .ZN(\sra_198/n266 ) );
  INV_X1 \sra_198/U223  ( .A(PR_1[8]), .ZN(\sra_198/n267 ) );
  INV_X1 \sra_198/U222  ( .A(PR_1[9]), .ZN(\sra_198/n268 ) );
  INV_X1 \sra_198/U221  ( .A(PR_1[10]), .ZN(\sra_198/n269 ) );
  INV_X1 \sra_198/U220  ( .A(PR_1[29]), .ZN(\sra_198/n288 ) );
  INV_X1 \sra_198/U219  ( .A(ct_1[4]), .ZN(\sra_198/n222 ) );
  INV_X1 \sra_198/U218  ( .A(PR_1[31]), .ZN(\sra_198/n260 ) );
  NAND2_X1 \sra_198/U217  ( .A1(ct_1[3]), .A2(PR_1[31]), .ZN(\sra_198/n163 )
         );
  INV_X1 \sra_198/U216  ( .A(ct_1[2]), .ZN(\sra_198/n245 ) );
  AOI22_X1 \sra_198/U215  ( .A1(PR_1[1]), .A2(\sra_198/n215 ), .B1(PR_1[0]), 
        .B2(\sra_198/n124 ), .ZN(\sra_198/n212 ) );
  INV_X1 \sra_198/U214  ( .A(ct_1[3]), .ZN(\sra_198/n243 ) );
  NAND2_X1 \sra_198/U213  ( .A1(ct_1[5]), .A2(PR_1[31]), .ZN(\sra_198/n112 )
         );
  NOR2_X1 \sra_198/U212  ( .A1(ct_1[4]), .A2(ct_1[5]), .ZN(\sra_198/n137 ) );
  NAND2_X1 \sra_198/U211  ( .A1(ct_1[2]), .A2(\sra_198/n243 ), .ZN(
        \sra_198/n146 ) );
  NOR2_X1 \sra_198/U210  ( .A1(\sra_198/n147 ), .A2(ct_1[4]), .ZN(
        \sra_198/n113 ) );
  NAND2_X1 \sra_198/U209  ( .A1(\sra_198/n196 ), .A2(ct_1[2]), .ZN(
        \sra_198/n74 ) );
  NAND2_X1 \sra_198/U208  ( .A1(PR_1[31]), .A2(\sra_198/n220 ), .ZN(
        \sra_198/n127 ) );
  AOI222_X1 \sra_198/U207  ( .A1(\sra_198/n88 ), .A2(\sra_198/n118 ), .B1(
        \sra_198/n86 ), .B2(\sra_198/n119 ), .C1(\sra_198/n110 ), .C2(
        \sra_198/n242 ), .ZN(\sra_198/n202 ) );
  AOI222_X1 \sra_198/U205  ( .A1(\sra_198/n82 ), .A2(\sra_198/n118 ), .B1(
        \sra_198/n78 ), .B2(\sra_198/n119 ), .C1(\sra_198/n106 ), .C2(
        \sra_198/n242 ), .ZN(\sra_198/n157 ) );
  AOI222_X1 \sra_198/U204  ( .A1(\sra_198/n99 ), .A2(\sra_198/n118 ), .B1(
        \sra_198/n102 ), .B2(\sra_198/n119 ), .C1(\sra_198/n101 ), .C2(
        \sra_198/n242 ), .ZN(\sra_198/n131 ) );
  AOI222_X1 \sra_198/U203  ( .A1(\sra_198/n92 ), .A2(\sra_198/n118 ), .B1(
        \sra_198/n95 ), .B2(\sra_198/n119 ), .C1(\sra_198/n94 ), .C2(
        \sra_198/n242 ), .ZN(\sra_198/n116 ) );
  INV_X1 \sra_198/U202  ( .A(ct_1[0]), .ZN(\sra_198/n259 ) );
  NOR2_X1 \sra_198/U201  ( .A1(ct_1[0]), .A2(ct_1[1]), .ZN(\sra_198/n124 ) );
  NOR2_X1 \sra_198/U200  ( .A1(\sra_198/n259 ), .A2(ct_1[1]), .ZN(
        \sra_198/n123 ) );
  OAI21_X1 \sra_198/U199  ( .B1(ct_1[5]), .B2(\sra_198/n199 ), .A(
        \sra_198/n112 ), .ZN(N264) );
  OAI21_X1 \sra_198/U198  ( .B1(ct_1[5]), .B2(\sra_198/n154 ), .A(
        \sra_198/n112 ), .ZN(N265) );
  OAI21_X1 \sra_198/U197  ( .B1(ct_1[5]), .B2(\sra_198/n128 ), .A(
        \sra_198/n112 ), .ZN(N266) );
  OAI21_X1 \sra_198/U196  ( .B1(ct_1[5]), .B2(\sra_198/n111 ), .A(
        \sra_198/n112 ), .ZN(N267) );
  INV_X1 \sra_198/U195  ( .A(PR_1[2]), .ZN(\sra_198/n261 ) );
  INV_X1 \sra_198/U194  ( .A(\sra_198/n201 ), .ZN(\sra_198/n226 ) );
  OAI221_X1 \sra_198/U193  ( .B1(\sra_198/n120 ), .B2(\sra_198/n261 ), .C1(
        \sra_198/n216 ), .C2(\sra_198/n262 ), .A(\sra_198/n212 ), .ZN(
        \sra_198/n200 ) );
  AOI21_X1 \sra_198/U192  ( .B1(\sra_198/n113 ), .B2(\sra_198/n200 ), .A(
        \sra_198/n226 ), .ZN(\sra_198/n199 ) );
  AOI22_X1 \sra_198/U191  ( .A1(PR_1[4]), .A2(\sra_198/n215 ), .B1(PR_1[3]), 
        .B2(\sra_198/n214 ), .ZN(\sra_198/n125 ) );
  INV_X1 \sra_198/U190  ( .A(\sra_198/n115 ), .ZN(\sra_198/n223 ) );
  OAI221_X1 \sra_198/U189  ( .B1(\sra_198/n120 ), .B2(\sra_198/n264 ), .C1(
        \sra_198/n216 ), .C2(\sra_198/n265 ), .A(\sra_198/n125 ), .ZN(
        \sra_198/n114 ) );
  AOI21_X1 \sra_198/U188  ( .B1(\sra_198/n113 ), .B2(\sra_198/n114 ), .A(
        \sra_198/n223 ), .ZN(\sra_198/n111 ) );
  AOI22_X1 \sra_198/U187  ( .A1(PR_1[2]), .A2(\sra_198/n123 ), .B1(PR_1[1]), 
        .B2(\sra_198/n214 ), .ZN(\sra_198/n161 ) );
  INV_X1 \sra_198/U186  ( .A(\sra_198/n156 ), .ZN(\sra_198/n225 ) );
  OAI221_X1 \sra_198/U185  ( .B1(\sra_198/n120 ), .B2(\sra_198/n262 ), .C1(
        \sra_198/n121 ), .C2(\sra_198/n263 ), .A(\sra_198/n161 ), .ZN(
        \sra_198/n155 ) );
  AOI21_X1 \sra_198/U184  ( .B1(\sra_198/n113 ), .B2(\sra_198/n155 ), .A(
        \sra_198/n225 ), .ZN(\sra_198/n154 ) );
  AOI22_X1 \sra_198/U183  ( .A1(PR_1[3]), .A2(\sra_198/n123 ), .B1(PR_1[2]), 
        .B2(\sra_198/n214 ), .ZN(\sra_198/n134 ) );
  INV_X1 \sra_198/U182  ( .A(\sra_198/n130 ), .ZN(\sra_198/n224 ) );
  OAI221_X1 \sra_198/U181  ( .B1(\sra_198/n120 ), .B2(\sra_198/n263 ), .C1(
        \sra_198/n121 ), .C2(\sra_198/n264 ), .A(\sra_198/n134 ), .ZN(
        \sra_198/n129 ) );
  AOI21_X1 \sra_198/U180  ( .B1(\sra_198/n113 ), .B2(\sra_198/n129 ), .A(
        \sra_198/n224 ), .ZN(\sra_198/n128 ) );
  NAND2_X1 \sra_198/U179  ( .A1(ct_1[1]), .A2(\sra_198/n259 ), .ZN(
        \sra_198/n120 ) );
  NAND2_X1 \sra_198/U178  ( .A1(ct_1[1]), .A2(ct_1[0]), .ZN(\sra_198/n121 ) );
  AOI22_X1 \sra_198/U177  ( .A1(PR_1[13]), .A2(\sra_198/n215 ), .B1(PR_1[12]), 
        .B2(\sra_198/n214 ), .ZN(\sra_198/n210 ) );
  OAI221_X1 \sra_198/U176  ( .B1(\sra_198/n120 ), .B2(\sra_198/n273 ), .C1(
        \sra_198/n216 ), .C2(\sra_198/n274 ), .A(\sra_198/n210 ), .ZN(
        \sra_198/n86 ) );
  AOI22_X1 \sra_198/U175  ( .A1(PR_1[9]), .A2(\sra_198/n215 ), .B1(PR_1[8]), 
        .B2(\sra_198/n124 ), .ZN(\sra_198/n211 ) );
  OAI221_X1 \sra_198/U174  ( .B1(\sra_198/n120 ), .B2(\sra_198/n269 ), .C1(
        \sra_198/n216 ), .C2(\sra_198/n270 ), .A(\sra_198/n211 ), .ZN(
        \sra_198/n88 ) );
  AOI22_X1 \sra_198/U173  ( .A1(PR_1[17]), .A2(\sra_198/n215 ), .B1(PR_1[16]), 
        .B2(\sra_198/n124 ), .ZN(\sra_198/n207 ) );
  OAI221_X1 \sra_198/U172  ( .B1(\sra_198/n120 ), .B2(\sra_198/n277 ), .C1(
        \sra_198/n216 ), .C2(\sra_198/n278 ), .A(\sra_198/n207 ), .ZN(
        \sra_198/n89 ) );
  AOI22_X1 \sra_198/U171  ( .A1(PR_1[18]), .A2(\sra_198/n123 ), .B1(PR_1[17]), 
        .B2(\sra_198/n124 ), .ZN(\sra_198/n177 ) );
  OAI221_X1 \sra_198/U170  ( .B1(\sra_198/n120 ), .B2(\sra_198/n278 ), .C1(
        \sra_198/n121 ), .C2(\sra_198/n279 ), .A(\sra_198/n177 ), .ZN(
        \sra_198/n83 ) );
  AOI22_X1 \sra_198/U169  ( .A1(PR_1[14]), .A2(\sra_198/n123 ), .B1(PR_1[13]), 
        .B2(\sra_198/n124 ), .ZN(\sra_198/n179 ) );
  OAI221_X1 \sra_198/U168  ( .B1(\sra_198/n217 ), .B2(\sra_198/n274 ), .C1(
        \sra_198/n121 ), .C2(\sra_198/n275 ), .A(\sra_198/n179 ), .ZN(
        \sra_198/n78 ) );
  AOI22_X1 \sra_198/U167  ( .A1(PR_1[19]), .A2(\sra_198/n215 ), .B1(PR_1[18]), 
        .B2(\sra_198/n214 ), .ZN(\sra_198/n195 ) );
  OAI221_X1 \sra_198/U166  ( .B1(\sra_198/n217 ), .B2(\sra_198/n279 ), .C1(
        \sra_198/n121 ), .C2(\sra_198/n280 ), .A(\sra_198/n195 ), .ZN(
        \sra_198/n166 ) );
  AOI22_X1 \sra_198/U165  ( .A1(PR_1[20]), .A2(\sra_198/n123 ), .B1(PR_1[19]), 
        .B2(\sra_198/n214 ), .ZN(\sra_198/n188 ) );
  OAI221_X1 \sra_198/U164  ( .B1(\sra_198/n217 ), .B2(\sra_198/n280 ), .C1(
        \sra_198/n121 ), .C2(\sra_198/n281 ), .A(\sra_198/n188 ), .ZN(
        \sra_198/n96 ) );
  AOI22_X1 \sra_198/U163  ( .A1(PR_1[22]), .A2(\sra_198/n123 ), .B1(PR_1[21]), 
        .B2(\sra_198/n124 ), .ZN(\sra_198/n178 ) );
  OAI221_X1 \sra_198/U162  ( .B1(\sra_198/n120 ), .B2(\sra_198/n282 ), .C1(
        \sra_198/n121 ), .C2(\sra_198/n283 ), .A(\sra_198/n178 ), .ZN(
        \sra_198/n152 ) );
  AOI22_X1 \sra_198/U161  ( .A1(PR_1[11]), .A2(\sra_198/n215 ), .B1(PR_1[10]), 
        .B2(\sra_198/n124 ), .ZN(\sra_198/n197 ) );
  OAI221_X1 \sra_198/U160  ( .B1(\sra_198/n217 ), .B2(\sra_198/n271 ), .C1(
        \sra_198/n121 ), .C2(\sra_198/n272 ), .A(\sra_198/n197 ), .ZN(
        \sra_198/n99 ) );
  AOI22_X1 \sra_198/U159  ( .A1(PR_1[15]), .A2(\sra_198/n215 ), .B1(PR_1[14]), 
        .B2(\sra_198/n214 ), .ZN(\sra_198/n194 ) );
  OAI221_X1 \sra_198/U158  ( .B1(\sra_198/n217 ), .B2(\sra_198/n275 ), .C1(
        \sra_198/n121 ), .C2(\sra_198/n276 ), .A(\sra_198/n194 ), .ZN(
        \sra_198/n102 ) );
  AOI22_X1 \sra_198/U157  ( .A1(PR_1[24]), .A2(\sra_198/n123 ), .B1(PR_1[23]), 
        .B2(\sra_198/n124 ), .ZN(\sra_198/n190 ) );
  OAI221_X1 \sra_198/U156  ( .B1(\sra_198/n217 ), .B2(\sra_198/n284 ), .C1(
        \sra_198/n121 ), .C2(\sra_198/n285 ), .A(\sra_198/n190 ), .ZN(
        \sra_198/n145 ) );
  AOI22_X1 \sra_198/U155  ( .A1(PR_1[12]), .A2(\sra_198/n215 ), .B1(PR_1[11]), 
        .B2(\sra_198/n214 ), .ZN(\sra_198/n189 ) );
  OAI221_X1 \sra_198/U154  ( .B1(\sra_198/n217 ), .B2(\sra_198/n272 ), .C1(
        \sra_198/n121 ), .C2(\sra_198/n273 ), .A(\sra_198/n189 ), .ZN(
        \sra_198/n92 ) );
  AOI22_X1 \sra_198/U153  ( .A1(PR_1[16]), .A2(\sra_198/n123 ), .B1(PR_1[15]), 
        .B2(\sra_198/n124 ), .ZN(\sra_198/n187 ) );
  OAI221_X1 \sra_198/U152  ( .B1(\sra_198/n217 ), .B2(\sra_198/n276 ), .C1(
        \sra_198/n121 ), .C2(\sra_198/n277 ), .A(\sra_198/n187 ), .ZN(
        \sra_198/n95 ) );
  AOI22_X1 \sra_198/U151  ( .A1(PR_1[25]), .A2(\sra_198/n215 ), .B1(PR_1[24]), 
        .B2(\sra_198/n214 ), .ZN(\sra_198/n205 ) );
  OAI221_X1 \sra_198/U150  ( .B1(\sra_198/n217 ), .B2(\sra_198/n285 ), .C1(
        \sra_198/n286 ), .C2(\sra_198/n216 ), .A(\sra_198/n205 ), .ZN(
        \sra_198/n143 ) );
  AOI22_X1 \sra_198/U149  ( .A1(PR_1[26]), .A2(\sra_198/n123 ), .B1(PR_1[25]), 
        .B2(\sra_198/n124 ), .ZN(\sra_198/n180 ) );
  OAI221_X1 \sra_198/U148  ( .B1(\sra_198/n217 ), .B2(\sra_198/n286 ), .C1(
        \sra_198/n121 ), .C2(\sra_198/n287 ), .A(\sra_198/n180 ), .ZN(
        \sra_198/n141 ) );
  AOI22_X1 \sra_198/U147  ( .A1(PR_1[27]), .A2(\sra_198/n215 ), .B1(PR_1[26]), 
        .B2(\sra_198/n214 ), .ZN(\sra_198/n193 ) );
  OAI221_X1 \sra_198/U146  ( .B1(\sra_198/n120 ), .B2(\sra_198/n287 ), .C1(
        \sra_198/n288 ), .C2(\sra_198/n216 ), .A(\sra_198/n193 ), .ZN(
        \sra_198/n164 ) );
  AOI22_X1 \sra_198/U145  ( .A1(PR_1[28]), .A2(\sra_198/n215 ), .B1(PR_1[27]), 
        .B2(\sra_198/n124 ), .ZN(\sra_198/n186 ) );
  OAI221_X1 \sra_198/U144  ( .B1(\sra_198/n288 ), .B2(\sra_198/n120 ), .C1(
        \sra_198/n289 ), .C2(\sra_198/n216 ), .A(\sra_198/n186 ), .ZN(
        \sra_198/n144 ) );
  AOI22_X1 \sra_198/U143  ( .A1(PR_1[29]), .A2(\sra_198/n215 ), .B1(PR_1[28]), 
        .B2(\sra_198/n214 ), .ZN(\sra_198/n206 ) );
  OAI221_X1 \sra_198/U141  ( .B1(\sra_198/n289 ), .B2(\sra_198/n120 ), .C1(
        \sra_198/n260 ), .C2(\sra_198/n216 ), .A(\sra_198/n206 ), .ZN(
        \sra_198/n142 ) );
  AOI22_X1 \sra_198/U140  ( .A1(PR_1[5]), .A2(\sra_198/n215 ), .B1(PR_1[4]), 
        .B2(\sra_198/n214 ), .ZN(\sra_198/n209 ) );
  OAI221_X1 \sra_198/U139  ( .B1(\sra_198/n120 ), .B2(\sra_198/n265 ), .C1(
        \sra_198/n216 ), .C2(\sra_198/n266 ), .A(\sra_198/n209 ), .ZN(
        \sra_198/n110 ) );
  AOI22_X1 \sra_198/U138  ( .A1(PR_1[8]), .A2(\sra_198/n215 ), .B1(PR_1[7]), 
        .B2(\sra_198/n214 ), .ZN(\sra_198/n122 ) );
  OAI221_X1 \sra_198/U137  ( .B1(\sra_198/n120 ), .B2(\sra_198/n268 ), .C1(
        \sra_198/n216 ), .C2(\sra_198/n269 ), .A(\sra_198/n122 ), .ZN(
        \sra_198/n94 ) );
  AOI22_X1 \sra_198/U136  ( .A1(PR_1[10]), .A2(\sra_198/n123 ), .B1(PR_1[9]), 
        .B2(\sra_198/n214 ), .ZN(\sra_198/n160 ) );
  OAI221_X1 \sra_198/U135  ( .B1(\sra_198/n120 ), .B2(\sra_198/n270 ), .C1(
        \sra_198/n121 ), .C2(\sra_198/n271 ), .A(\sra_198/n160 ), .ZN(
        \sra_198/n82 ) );
  AOI22_X1 \sra_198/U134  ( .A1(PR_1[6]), .A2(\sra_198/n215 ), .B1(PR_1[5]), 
        .B2(\sra_198/n214 ), .ZN(\sra_198/n159 ) );
  OAI221_X1 \sra_198/U133  ( .B1(\sra_198/n120 ), .B2(\sra_198/n266 ), .C1(
        \sra_198/n121 ), .C2(\sra_198/n267 ), .A(\sra_198/n159 ), .ZN(
        \sra_198/n106 ) );
  AOI22_X1 \sra_198/U132  ( .A1(PR_1[7]), .A2(\sra_198/n215 ), .B1(PR_1[6]), 
        .B2(\sra_198/n214 ), .ZN(\sra_198/n133 ) );
  OAI221_X1 \sra_198/U131  ( .B1(\sra_198/n120 ), .B2(\sra_198/n267 ), .C1(
        \sra_198/n216 ), .C2(\sra_198/n268 ), .A(\sra_198/n133 ), .ZN(
        \sra_198/n101 ) );
  OAI211_X1 \sra_198/U130  ( .C1(\sra_198/n248 ), .C2(\sra_198/n74 ), .A(
        \sra_198/n107 ), .B(\sra_198/n108 ), .ZN(N268) );
  OAI211_X1 \sra_198/U129  ( .C1(\sra_198/n249 ), .C2(\sra_198/n74 ), .A(
        \sra_198/n103 ), .B(\sra_198/n104 ), .ZN(N269) );
  OAI211_X1 \sra_198/U128  ( .C1(\sra_198/n256 ), .C2(\sra_198/n74 ), .A(
        \sra_198/n97 ), .B(\sra_198/n98 ), .ZN(N270) );
  OAI211_X1 \sra_198/U127  ( .C1(\sra_198/n253 ), .C2(\sra_198/n74 ), .A(
        \sra_198/n90 ), .B(\sra_198/n91 ), .ZN(N271) );
  OAI211_X1 \sra_198/U126  ( .C1(\sra_198/n247 ), .C2(\sra_198/n74 ), .A(
        \sra_198/n84 ), .B(\sra_198/n85 ), .ZN(N272) );
  OAI211_X1 \sra_198/U125  ( .C1(\sra_198/n250 ), .C2(\sra_198/n74 ), .A(
        \sra_198/n75 ), .B(\sra_198/n76 ), .ZN(N273) );
  OAI211_X1 \sra_198/U124  ( .C1(\sra_198/n257 ), .C2(\sra_198/n74 ), .A(
        \sra_198/n191 ), .B(\sra_198/n192 ), .ZN(N274) );
  OAI211_X1 \sra_198/U123  ( .C1(\sra_198/n254 ), .C2(\sra_198/n74 ), .A(
        \sra_198/n184 ), .B(\sra_198/n185 ), .ZN(N275) );
  OAI211_X1 \sra_198/U122  ( .C1(\sra_198/n258 ), .C2(\sra_198/n74 ), .A(
        \sra_198/n181 ), .B(\sra_198/n182 ), .ZN(N276) );
  OAI211_X1 \sra_198/U121  ( .C1(\sra_198/n251 ), .C2(\sra_198/n74 ), .A(
        \sra_198/n175 ), .B(\sra_198/n176 ), .ZN(N277) );
  OAI211_X1 \sra_198/U120  ( .C1(\sra_198/n255 ), .C2(\sra_198/n74 ), .A(
        \sra_198/n171 ), .B(\sra_198/n172 ), .ZN(N278) );
  OAI221_X1 \sra_198/U119  ( .B1(\sra_198/n254 ), .B2(\sra_198/n169 ), .C1(
        \sra_198/n252 ), .C2(\sra_198/n74 ), .A(\sra_198/n170 ), .ZN(N279) );
  OAI21_X1 \sra_198/U118  ( .B1(\sra_198/n239 ), .B2(\sra_198/n220 ), .A(
        \sra_198/n127 ), .ZN(N280) );
  OAI21_X1 \sra_198/U117  ( .B1(\sra_198/n158 ), .B2(\sra_198/n220 ), .A(
        \sra_198/n127 ), .ZN(N281) );
  OAI21_X1 \sra_198/U116  ( .B1(\sra_198/n132 ), .B2(\sra_198/n220 ), .A(
        \sra_198/n127 ), .ZN(N282) );
  OAI21_X1 \sra_198/U114  ( .B1(\sra_198/n117 ), .B2(\sra_198/n220 ), .A(
        \sra_198/n127 ), .ZN(N283) );
  OAI21_X1 \sra_198/U113  ( .B1(\sra_198/n238 ), .B2(\sra_198/n220 ), .A(
        \sra_198/n127 ), .ZN(N284) );
  OAI21_X1 \sra_198/U112  ( .B1(\sra_198/n237 ), .B2(\sra_198/n220 ), .A(
        \sra_198/n127 ), .ZN(N285) );
  OAI21_X1 \sra_198/U111  ( .B1(\sra_198/n236 ), .B2(\sra_198/n220 ), .A(
        \sra_198/n127 ), .ZN(N286) );
  OAI21_X1 \sra_198/U110  ( .B1(\sra_198/n93 ), .B2(\sra_198/n220 ), .A(
        \sra_198/n127 ), .ZN(N287) );
  OAI21_X1 \sra_198/U109  ( .B1(\sra_198/n87 ), .B2(\sra_198/n220 ), .A(
        \sra_198/n127 ), .ZN(N288) );
  OAI21_X1 \sra_198/U108  ( .B1(\sra_198/n80 ), .B2(\sra_198/n220 ), .A(
        \sra_198/n127 ), .ZN(N289) );
  OAI21_X1 \sra_198/U107  ( .B1(\sra_198/n140 ), .B2(\sra_198/n220 ), .A(
        \sra_198/n127 ), .ZN(N290) );
  OAI21_X1 \sra_198/U105  ( .B1(\sra_198/n139 ), .B2(\sra_198/n220 ), .A(
        \sra_198/n127 ), .ZN(N291) );
  OAI21_X1 \sra_198/U104  ( .B1(\sra_198/n138 ), .B2(\sra_198/n220 ), .A(
        \sra_198/n127 ), .ZN(N292) );
  INV_X1 \sra_198/U103  ( .A(\sra_198/n135 ), .ZN(N293) );
  OAI21_X1 \sra_198/U102  ( .B1(\sra_198/n126 ), .B2(\sra_198/n220 ), .A(
        \sra_198/n127 ), .ZN(N294) );
  AOI22_X1 \sra_198/U101  ( .A1(PR_1[21]), .A2(\sra_198/n215 ), .B1(PR_1[20]), 
        .B2(\sra_198/n214 ), .ZN(\sra_198/n208 ) );
  OAI221_X1 \sra_198/U100  ( .B1(\sra_198/n217 ), .B2(\sra_198/n281 ), .C1(
        \sra_198/n121 ), .C2(\sra_198/n282 ), .A(\sra_198/n208 ), .ZN(
        \sra_198/n183 ) );
  AOI22_X1 \sra_198/U99  ( .A1(PR_1[23]), .A2(\sra_198/n215 ), .B1(PR_1[22]), 
        .B2(\sra_198/n214 ), .ZN(\sra_198/n198 ) );
  OAI221_X1 \sra_198/U98  ( .B1(\sra_198/n217 ), .B2(\sra_198/n283 ), .C1(
        \sra_198/n216 ), .C2(\sra_198/n284 ), .A(\sra_198/n198 ), .ZN(
        \sra_198/n174 ) );
  AOI222_X1 \sra_198/U97  ( .A1(\sra_198/n214 ), .A2(PR_1[29]), .B1(
        \sra_198/n123 ), .B2(PR_1[30]), .C1(PR_1[31]), .C2(ct_1[1]), .ZN(
        \sra_198/n168 ) );
  INV_X1 \sra_198/U96  ( .A(\sra_198/n126 ), .ZN(\sra_198/n229 ) );
  AOI221_X1 \sra_198/U95  ( .B1(\sra_198/n77 ), .B2(\sra_198/n166 ), .C1(
        \sra_198/n79 ), .C2(\sra_198/n229 ), .A(\sra_198/n221 ), .ZN(
        \sra_198/n172 ) );
  INV_X1 \sra_198/U94  ( .A(\sra_198/n83 ), .ZN(\sra_198/n249 ) );
  INV_X1 \sra_198/U93  ( .A(\sra_198/n144 ), .ZN(\sra_198/n252 ) );
  NAND2_X1 \sra_198/U92  ( .A1(\sra_198/n196 ), .A2(\sra_198/n245 ), .ZN(
        \sra_198/n169 ) );
  INV_X1 \sra_198/U91  ( .A(\sra_198/n96 ), .ZN(\sra_198/n253 ) );
  INV_X1 \sra_198/U90  ( .A(\sra_198/n145 ), .ZN(\sra_198/n254 ) );
  INV_X1 \sra_198/U89  ( .A(\sra_198/n127 ), .ZN(\sra_198/n219 ) );
  INV_X1 \sra_198/U88  ( .A(\sra_198/n163 ), .ZN(\sra_198/n244 ) );
  AOI21_X1 \sra_198/U87  ( .B1(\sra_198/n136 ), .B2(\sra_198/n137 ), .A(
        \sra_198/n219 ), .ZN(\sra_198/n135 ) );
  NOR2_X1 \sra_198/U86  ( .A1(\sra_198/n220 ), .A2(\sra_198/n243 ), .ZN(
        \sra_198/n196 ) );
  INV_X1 \sra_198/U85  ( .A(\sra_198/n173 ), .ZN(\sra_198/n228 ) );
  OAI21_X1 \sra_198/U84  ( .B1(\sra_198/n168 ), .B2(\sra_198/n147 ), .A(
        \sra_198/n228 ), .ZN(\sra_198/n136 ) );
  AOI21_X1 \sra_198/U83  ( .B1(\sra_198/n149 ), .B2(\sra_198/n235 ), .A(
        \sra_198/n173 ), .ZN(\sra_198/n126 ) );
  AOI22_X1 \sra_198/U82  ( .A1(\sra_198/n81 ), .A2(\sra_198/n110 ), .B1(
        \sra_198/n218 ), .B2(\sra_198/n86 ), .ZN(\sra_198/n107 ) );
  AOI22_X1 \sra_198/U81  ( .A1(\sra_198/n81 ), .A2(\sra_198/n106 ), .B1(
        \sra_198/n218 ), .B2(\sra_198/n78 ), .ZN(\sra_198/n103 ) );
  AOI22_X1 \sra_198/U80  ( .A1(\sra_198/n81 ), .A2(\sra_198/n101 ), .B1(
        \sra_198/n218 ), .B2(\sra_198/n102 ), .ZN(\sra_198/n97 ) );
  AOI22_X1 \sra_198/U79  ( .A1(\sra_198/n81 ), .A2(\sra_198/n94 ), .B1(
        \sra_198/n218 ), .B2(\sra_198/n95 ), .ZN(\sra_198/n90 ) );
  AOI22_X1 \sra_198/U78  ( .A1(\sra_198/n81 ), .A2(\sra_198/n88 ), .B1(
        \sra_198/n218 ), .B2(\sra_198/n89 ), .ZN(\sra_198/n84 ) );
  AOI22_X1 \sra_198/U77  ( .A1(\sra_198/n81 ), .A2(\sra_198/n82 ), .B1(
        \sra_198/n218 ), .B2(\sra_198/n83 ), .ZN(\sra_198/n75 ) );
  AOI22_X1 \sra_198/U76  ( .A1(\sra_198/n81 ), .A2(\sra_198/n99 ), .B1(
        \sra_198/n218 ), .B2(\sra_198/n166 ), .ZN(\sra_198/n191 ) );
  AOI22_X1 \sra_198/U75  ( .A1(\sra_198/n81 ), .A2(\sra_198/n92 ), .B1(
        \sra_198/n218 ), .B2(\sra_198/n96 ), .ZN(\sra_198/n184 ) );
  AOI22_X1 \sra_198/U74  ( .A1(\sra_198/n81 ), .A2(\sra_198/n86 ), .B1(
        \sra_198/n218 ), .B2(\sra_198/n183 ), .ZN(\sra_198/n181 ) );
  AOI22_X1 \sra_198/U73  ( .A1(\sra_198/n81 ), .A2(\sra_198/n78 ), .B1(
        \sra_198/n218 ), .B2(\sra_198/n152 ), .ZN(\sra_198/n175 ) );
  AOI22_X1 \sra_198/U72  ( .A1(\sra_198/n81 ), .A2(\sra_198/n102 ), .B1(
        \sra_198/n218 ), .B2(\sra_198/n174 ), .ZN(\sra_198/n171 ) );
  NOR2_X1 \sra_198/U71  ( .A1(\sra_198/n163 ), .A2(\sra_198/n245 ), .ZN(
        \sra_198/n150 ) );
  NOR2_X1 \sra_198/U70  ( .A1(\sra_198/n260 ), .A2(\sra_198/n235 ), .ZN(
        \sra_198/n173 ) );
  AOI221_X1 \sra_198/U69  ( .B1(\sra_198/n77 ), .B2(\sra_198/n83 ), .C1(
        \sra_198/n79 ), .C2(\sra_198/n136 ), .A(\sra_198/n221 ), .ZN(
        \sra_198/n176 ) );
  INV_X1 \sra_198/U68  ( .A(\sra_198/n137 ), .ZN(\sra_198/n220 ) );
  AOI221_X1 \sra_198/U67  ( .B1(\sra_198/n81 ), .B2(\sra_198/n95 ), .C1(
        \sra_198/n77 ), .C2(\sra_198/n96 ), .A(\sra_198/n219 ), .ZN(
        \sra_198/n170 ) );
  NAND2_X1 \sra_198/U66  ( .A1(\sra_198/n245 ), .A2(\sra_198/n243 ), .ZN(
        \sra_198/n147 ) );
  INV_X1 \sra_198/U65  ( .A(\sra_198/n146 ), .ZN(\sra_198/n242 ) );
  INV_X1 \sra_198/U64  ( .A(\sra_198/n112 ), .ZN(\sra_198/n221 ) );
  NOR2_X1 \sra_198/U63  ( .A1(\sra_198/n245 ), .A2(\sra_198/n243 ), .ZN(
        \sra_198/n119 ) );
  INV_X1 \sra_198/U62  ( .A(\sra_198/n139 ), .ZN(\sra_198/n231 ) );
  AOI221_X1 \sra_198/U61  ( .B1(\sra_198/n77 ), .B2(\sra_198/n95 ), .C1(
        \sra_198/n79 ), .C2(\sra_198/n231 ), .A(\sra_198/n221 ), .ZN(
        \sra_198/n185 ) );
  INV_X1 \sra_198/U60  ( .A(\sra_198/n138 ), .ZN(\sra_198/n230 ) );
  AOI221_X1 \sra_198/U59  ( .B1(\sra_198/n77 ), .B2(\sra_198/n89 ), .C1(
        \sra_198/n79 ), .C2(\sra_198/n230 ), .A(\sra_198/n221 ), .ZN(
        \sra_198/n182 ) );
  INV_X1 \sra_198/U58  ( .A(\sra_198/n89 ), .ZN(\sra_198/n248 ) );
  INV_X1 \sra_198/U57  ( .A(\sra_198/n152 ), .ZN(\sra_198/n250 ) );
  INV_X1 \sra_198/U56  ( .A(\sra_198/n164 ), .ZN(\sra_198/n255 ) );
  INV_X1 \sra_198/U55  ( .A(\sra_198/n166 ), .ZN(\sra_198/n256 ) );
  INV_X1 \sra_198/U54  ( .A(\sra_198/n143 ), .ZN(\sra_198/n258 ) );
  INV_X1 \sra_198/U53  ( .A(\sra_198/n141 ), .ZN(\sra_198/n251 ) );
  INV_X1 \sra_198/U52  ( .A(\sra_198/n174 ), .ZN(\sra_198/n257 ) );
  INV_X1 \sra_198/U51  ( .A(\sra_198/n183 ), .ZN(\sra_198/n247 ) );
  INV_X1 \sra_198/U50  ( .A(\sra_198/n168 ), .ZN(\sra_198/n246 ) );
  BUF_X1 \sra_198/U49  ( .A(\sra_198/n124 ), .Z(\sra_198/n214 ) );
  AOI21_X1 \sra_198/U48  ( .B1(\sra_198/n118 ), .B2(\sra_198/n142 ), .A(
        \sra_198/n150 ), .ZN(\sra_198/n153 ) );
  OAI221_X1 \sra_198/U47  ( .B1(\sra_198/n258 ), .B2(\sra_198/n146 ), .C1(
        \sra_198/n247 ), .C2(\sra_198/n147 ), .A(\sra_198/n153 ), .ZN(
        \sra_198/n109 ) );
  AOI22_X1 \sra_198/U46  ( .A1(\sra_198/n119 ), .A2(\sra_198/n142 ), .B1(
        \sra_198/n118 ), .B2(\sra_198/n143 ), .ZN(\sra_198/n204 ) );
  OAI221_X1 \sra_198/U45  ( .B1(\sra_198/n247 ), .B2(\sra_198/n146 ), .C1(
        \sra_198/n248 ), .C2(\sra_198/n147 ), .A(\sra_198/n204 ), .ZN(
        \sra_198/n203 ) );
  INV_X1 \sra_198/U44  ( .A(\sra_198/n203 ), .ZN(\sra_198/n239 ) );
  BUF_X1 \sra_198/U43  ( .A(\sra_198/n121 ), .Z(\sra_198/n216 ) );
  BUF_X1 \sra_198/U42  ( .A(\sra_198/n120 ), .Z(\sra_198/n217 ) );
  BUF_X1 \sra_198/U41  ( .A(\sra_198/n123 ), .Z(\sra_198/n215 ) );
  AOI21_X1 \sra_198/U40  ( .B1(\sra_198/n144 ), .B2(\sra_198/n235 ), .A(
        \sra_198/n173 ), .ZN(\sra_198/n139 ) );
  AOI21_X1 \sra_198/U39  ( .B1(\sra_198/n142 ), .B2(\sra_198/n235 ), .A(
        \sra_198/n173 ), .ZN(\sra_198/n138 ) );
  AOI221_X1 \sra_198/U38  ( .B1(\sra_198/n77 ), .B2(\sra_198/n88 ), .C1(
        \sra_198/n79 ), .C2(\sra_198/n109 ), .A(\sra_198/n221 ), .ZN(
        \sra_198/n108 ) );
  AOI221_X1 \sra_198/U37  ( .B1(\sra_198/n77 ), .B2(\sra_198/n82 ), .C1(
        \sra_198/n79 ), .C2(\sra_198/n105 ), .A(\sra_198/n221 ), .ZN(
        \sra_198/n104 ) );
  AOI221_X1 \sra_198/U36  ( .B1(\sra_198/n77 ), .B2(\sra_198/n99 ), .C1(
        \sra_198/n79 ), .C2(\sra_198/n100 ), .A(\sra_198/n221 ), .ZN(
        \sra_198/n98 ) );
  INV_X1 \sra_198/U35  ( .A(\sra_198/n93 ), .ZN(\sra_198/n232 ) );
  AOI221_X1 \sra_198/U34  ( .B1(\sra_198/n77 ), .B2(\sra_198/n92 ), .C1(
        \sra_198/n79 ), .C2(\sra_198/n232 ), .A(\sra_198/n221 ), .ZN(
        \sra_198/n91 ) );
  INV_X1 \sra_198/U33  ( .A(\sra_198/n87 ), .ZN(\sra_198/n233 ) );
  AOI221_X1 \sra_198/U32  ( .B1(\sra_198/n77 ), .B2(\sra_198/n86 ), .C1(
        \sra_198/n79 ), .C2(\sra_198/n233 ), .A(\sra_198/n221 ), .ZN(
        \sra_198/n85 ) );
  INV_X1 \sra_198/U31  ( .A(\sra_198/n80 ), .ZN(\sra_198/n234 ) );
  AOI221_X1 \sra_198/U30  ( .B1(\sra_198/n77 ), .B2(\sra_198/n78 ), .C1(
        \sra_198/n79 ), .C2(\sra_198/n234 ), .A(\sra_198/n221 ), .ZN(
        \sra_198/n76 ) );
  INV_X1 \sra_198/U29  ( .A(\sra_198/n140 ), .ZN(\sra_198/n227 ) );
  AOI221_X1 \sra_198/U28  ( .B1(\sra_198/n77 ), .B2(\sra_198/n102 ), .C1(
        \sra_198/n79 ), .C2(\sra_198/n227 ), .A(\sra_198/n221 ), .ZN(
        \sra_198/n192 ) );
  AOI21_X1 \sra_198/U27  ( .B1(\sra_198/n118 ), .B2(\sra_198/n246 ), .A(
        \sra_198/n150 ), .ZN(\sra_198/n151 ) );
  OAI221_X1 \sra_198/U26  ( .B1(\sra_198/n251 ), .B2(\sra_198/n146 ), .C1(
        \sra_198/n250 ), .C2(\sra_198/n147 ), .A(\sra_198/n151 ), .ZN(
        \sra_198/n105 ) );
  AOI21_X1 \sra_198/U25  ( .B1(\sra_198/n118 ), .B2(\sra_198/n149 ), .A(
        \sra_198/n150 ), .ZN(\sra_198/n148 ) );
  OAI221_X1 \sra_198/U24  ( .B1(\sra_198/n255 ), .B2(\sra_198/n146 ), .C1(
        \sra_198/n257 ), .C2(\sra_198/n147 ), .A(\sra_198/n148 ), .ZN(
        \sra_198/n100 ) );
  OAI22_X1 \sra_198/U23  ( .A1(\sra_198/n146 ), .A2(\sra_198/n257 ), .B1(
        \sra_198/n147 ), .B2(\sra_198/n256 ), .ZN(\sra_198/n165 ) );
  AOI221_X1 \sra_198/U22  ( .B1(\sra_198/n149 ), .B2(\sra_198/n119 ), .C1(
        \sra_198/n164 ), .C2(\sra_198/n118 ), .A(\sra_198/n165 ), .ZN(
        \sra_198/n132 ) );
  AOI22_X1 \sra_198/U21  ( .A1(\sra_198/n119 ), .A2(\sra_198/n246 ), .B1(
        \sra_198/n118 ), .B2(\sra_198/n141 ), .ZN(\sra_198/n167 ) );
  INV_X1 \sra_198/U20  ( .A(\sra_198/n167 ), .ZN(\sra_198/n241 ) );
  AOI221_X1 \sra_198/U19  ( .B1(\sra_198/n152 ), .B2(\sra_198/n242 ), .C1(
        \sra_198/n83 ), .C2(\sra_198/n235 ), .A(\sra_198/n241 ), .ZN(
        \sra_198/n158 ) );
  AOI21_X1 \sra_198/U18  ( .B1(\sra_198/n118 ), .B2(\sra_198/n144 ), .A(
        \sra_198/n150 ), .ZN(\sra_198/n162 ) );
  INV_X1 \sra_198/U17  ( .A(\sra_198/n162 ), .ZN(\sra_198/n240 ) );
  AOI221_X1 \sra_198/U16  ( .B1(\sra_198/n145 ), .B2(\sra_198/n242 ), .C1(
        \sra_198/n96 ), .C2(\sra_198/n235 ), .A(\sra_198/n240 ), .ZN(
        \sra_198/n117 ) );
  AOI221_X1 \sra_198/U15  ( .B1(\sra_198/n144 ), .B2(\sra_198/n242 ), .C1(
        \sra_198/n145 ), .C2(\sra_198/n235 ), .A(\sra_198/n244 ), .ZN(
        \sra_198/n93 ) );
  AOI221_X1 \sra_198/U14  ( .B1(\sra_198/n142 ), .B2(\sra_198/n242 ), .C1(
        \sra_198/n143 ), .C2(\sra_198/n235 ), .A(\sra_198/n244 ), .ZN(
        \sra_198/n87 ) );
  AOI221_X1 \sra_198/U13  ( .B1(\sra_198/n246 ), .B2(\sra_198/n242 ), .C1(
        \sra_198/n141 ), .C2(\sra_198/n235 ), .A(\sra_198/n244 ), .ZN(
        \sra_198/n80 ) );
  AOI221_X1 \sra_198/U12  ( .B1(\sra_198/n149 ), .B2(\sra_198/n242 ), .C1(
        \sra_198/n164 ), .C2(\sra_198/n235 ), .A(\sra_198/n244 ), .ZN(
        \sra_198/n140 ) );
  INV_X1 \sra_198/U11  ( .A(\sra_198/n105 ), .ZN(\sra_198/n237 ) );
  INV_X1 \sra_198/U10  ( .A(\sra_198/n100 ), .ZN(\sra_198/n236 ) );
  INV_X1 \sra_198/U9  ( .A(\sra_198/n169 ), .ZN(\sra_198/n218 ) );
  INV_X1 \sra_198/U8  ( .A(\sra_198/n147 ), .ZN(\sra_198/n235 ) );
  NOR2_X1 \sra_198/U7  ( .A1(\sra_198/n220 ), .A2(\sra_198/n147 ), .ZN(
        \sra_198/n81 ) );
  INV_X1 \sra_198/U6  ( .A(\sra_198/n109 ), .ZN(\sra_198/n238 ) );
  NOR2_X1 \sra_198/U5  ( .A1(\sra_198/n243 ), .A2(ct_1[2]), .ZN(\sra_198/n118 ) );
  NOR2_X1 \sra_198/U4  ( .A1(\sra_198/n222 ), .A2(ct_1[5]), .ZN(\sra_198/n79 )
         );
  NOR2_X1 \sra_198/U3  ( .A1(\sra_198/n220 ), .A2(\sra_198/n146 ), .ZN(
        \sra_198/n77 ) );
  MUX2_X1 \sra_198/U226  ( .A(\sra_198/n202 ), .B(\sra_198/n239 ), .S(ct_1[4]), 
        .Z(\sra_198/n201 ) );
  MUX2_X1 \sra_198/U206  ( .A(PR_1[31]), .B(PR_1[30]), .S(\sra_198/n214 ), .Z(
        \sra_198/n149 ) );
  MUX2_X1 \sra_198/U142  ( .A(\sra_198/n157 ), .B(\sra_198/n158 ), .S(ct_1[4]), 
        .Z(\sra_198/n156 ) );
  MUX2_X1 \sra_198/U115  ( .A(\sra_198/n131 ), .B(\sra_198/n132 ), .S(ct_1[4]), 
        .Z(\sra_198/n130 ) );
  MUX2_X1 \sra_198/U106  ( .A(\sra_198/n116 ), .B(\sra_198/n117 ), .S(ct_1[4]), 
        .Z(\sra_198/n115 ) );
  INV_X1 \add_35/U6  ( .A(q[0]), .ZN(qp1[0]) );
  XOR2_X1 \add_35/U5  ( .A(q[1]), .B(q[0]), .Z(qp1[1]) );
  XNOR2_X1 \add_35/U4  ( .A(\add_35/carry[30] ), .B(\add_35/n3 ), .ZN(qp1[30])
         );
  AND4_X1 \add_35/U3  ( .A1(q[16]), .A2(\add_35/carry[16] ), .A3(q[17]), .A4(
        q[18]), .ZN(\add_35/carry[19] ) );
  AND2_X1 \add_35/U2  ( .A1(q[1]), .A2(q[0]), .ZN(\add_35/n2 ) );
  INV_X1 \add_35/U1  ( .A(q[30]), .ZN(\add_35/n3 ) );
  HA_X1 \add_35/U1_1_2  ( .A(q[2]), .B(\add_35/n2 ), .CO(\add_35/carry[3] ), 
        .S(qp1[2]) );
  HA_X1 \add_35/U1_1_3  ( .A(\add_35/carry[3] ), .B(q[3]), .CO(
        \add_35/carry[4] ), .S(qp1[3]) );
  HA_X1 \add_35/U1_1_4  ( .A(\add_35/carry[4] ), .B(q[4]), .CO(
        \add_35/carry[5] ), .S(qp1[4]) );
  HA_X1 \add_35/U1_1_5  ( .A(\add_35/carry[5] ), .B(q[5]), .CO(
        \add_35/carry[6] ), .S(qp1[5]) );
  HA_X1 \add_35/U1_1_6  ( .A(\add_35/carry[6] ), .B(q[6]), .CO(
        \add_35/carry[7] ), .S(qp1[6]) );
  HA_X1 \add_35/U1_1_7  ( .A(\add_35/carry[7] ), .B(q[7]), .CO(
        \add_35/carry[8] ), .S(qp1[7]) );
  HA_X1 \add_35/U1_1_8  ( .A(\add_35/carry[8] ), .B(q[8]), .CO(
        \add_35/carry[9] ), .S(qp1[8]) );
  HA_X1 \add_35/U1_1_9  ( .A(\add_35/carry[9] ), .B(q[9]), .CO(
        \add_35/carry[10] ), .S(qp1[9]) );
  HA_X1 \add_35/U1_1_10  ( .A(\add_35/carry[10] ), .B(q[10]), .CO(
        \add_35/carry[11] ), .S(qp1[10]) );
  HA_X1 \add_35/U1_1_11  ( .A(\add_35/carry[11] ), .B(q[11]), .CO(
        \add_35/carry[12] ), .S(qp1[11]) );
  HA_X1 \add_35/U1_1_12  ( .A(q[12]), .B(\add_35/carry[12] ), .CO(
        \add_35/carry[13] ), .S(qp1[12]) );
  HA_X1 \add_35/U1_1_13  ( .A(\add_35/carry[13] ), .B(q[13]), .CO(
        \add_35/carry[14] ), .S(qp1[13]) );
  HA_X1 \add_35/U1_1_14  ( .A(\add_35/carry[14] ), .B(q[14]), .CO(
        \add_35/carry[15] ), .S(qp1[14]) );
  HA_X1 \add_35/U1_1_15  ( .A(\add_35/carry[15] ), .B(q[15]), .CO(
        \add_35/carry[16] ), .S(qp1[15]) );
  HA_X1 \add_35/U1_1_16  ( .A(q[16]), .B(\add_35/carry[16] ), .CO(
        \add_35/carry[17] ), .S(qp1[16]) );
  HA_X1 \add_35/U1_1_17  ( .A(\add_35/carry[17] ), .B(q[17]), .CO(
        \add_35/carry[18] ), .S(qp1[17]) );
  HA_X1 \add_35/U1_1_18  ( .A(\add_35/carry[18] ), .B(q[18]), .CO(), .S(
        qp1[18]) );
  HA_X1 \add_35/U1_1_19  ( .A(q[19]), .B(\add_35/carry[19] ), .CO(
        \add_35/carry[20] ), .S(qp1[19]) );
  HA_X1 \add_35/U1_1_20  ( .A(\add_35/carry[20] ), .B(q[20]), .CO(
        \add_35/carry[21] ), .S(qp1[20]) );
  HA_X1 \add_35/U1_1_21  ( .A(\add_35/carry[21] ), .B(q[21]), .CO(
        \add_35/carry[22] ), .S(qp1[21]) );
  HA_X1 \add_35/U1_1_22  ( .A(\add_35/carry[22] ), .B(q[22]), .CO(
        \add_35/carry[23] ), .S(qp1[22]) );
  HA_X1 \add_35/U1_1_23  ( .A(\add_35/carry[23] ), .B(q[23]), .CO(
        \add_35/carry[24] ), .S(qp1[23]) );
  HA_X1 \add_35/U1_1_24  ( .A(\add_35/carry[24] ), .B(q[24]), .CO(
        \add_35/carry[25] ), .S(qp1[24]) );
  HA_X1 \add_35/U1_1_25  ( .A(\add_35/carry[25] ), .B(q[25]), .CO(
        \add_35/carry[26] ), .S(qp1[25]) );
  HA_X1 \add_35/U1_1_26  ( .A(\add_35/carry[26] ), .B(q[26]), .CO(
        \add_35/carry[27] ), .S(qp1[26]) );
  HA_X1 \add_35/U1_1_27  ( .A(\add_35/carry[27] ), .B(q[27]), .CO(
        \add_35/carry[28] ), .S(qp1[27]) );
  HA_X1 \add_35/U1_1_28  ( .A(\add_35/carry[28] ), .B(q[28]), .CO(
        \add_35/carry[29] ), .S(qp1[28]) );
  HA_X1 \add_35/U1_1_29  ( .A(\add_35/carry[29] ), .B(q[29]), .CO(
        \add_35/carry[30] ), .S(qp1[29]) );
  INV_X1 \add_34/U11  ( .A(\add_34/n6 ), .ZN(nqp1[0]) );
  CLKBUF_X1 \add_34/U10  ( .A(n2931), .Z(\add_34/n6 ) );
  XNOR2_X1 \add_34/U9  ( .A(\add_34/carry[30] ), .B(\add_34/n5 ), .ZN(nqp1[30]) );
  INV_X1 \add_34/U8  ( .A(nq[30]), .ZN(\add_34/n5 ) );
  XOR2_X1 \add_34/U7  ( .A(n2930), .B(\add_34/n6 ), .Z(nqp1[1]) );
  AND2_X1 \add_34/U6  ( .A1(n2930), .A2(n2931), .ZN(\add_34/n4 ) );
  AND4_X1 \add_34/U5  ( .A1(\add_34/carry[26] ), .A2(nq[26]), .A3(nq[27]), 
        .A4(nq[28]), .ZN(\add_34/carry[29] ) );
  INV_X1 \add_34/U4  ( .A(\add_34/n3 ), .ZN(nqp1[28]) );
  XNOR2_X1 \add_34/U3  ( .A(\add_34/carry[28] ), .B(nq[28]), .ZN(\add_34/n3 )
         );
  AND3_X1 \add_34/U2  ( .A1(\add_34/carry[24] ), .A2(nq[24]), .A3(nq[25]), 
        .ZN(\add_34/carry[26] ) );
  CLKBUF_X1 \add_34/U1  ( .A(\add_34/carry[24] ), .Z(\add_34/n2 ) );
  HA_X1 \add_34/U1_1_2  ( .A(\add_34/n4 ), .B(nq[2]), .CO(\add_34/carry[3] ), 
        .S(nqp1[2]) );
  HA_X1 \add_34/U1_1_3  ( .A(\add_34/carry[3] ), .B(nq[3]), .CO(
        \add_34/carry[4] ), .S(nqp1[3]) );
  HA_X1 \add_34/U1_1_4  ( .A(\add_34/carry[4] ), .B(nq[4]), .CO(
        \add_34/carry[5] ), .S(nqp1[4]) );
  HA_X1 \add_34/U1_1_5  ( .A(\add_34/carry[5] ), .B(nq[5]), .CO(
        \add_34/carry[6] ), .S(nqp1[5]) );
  HA_X1 \add_34/U1_1_6  ( .A(\add_34/carry[6] ), .B(nq[6]), .CO(
        \add_34/carry[7] ), .S(nqp1[6]) );
  HA_X1 \add_34/U1_1_7  ( .A(\add_34/carry[7] ), .B(nq[7]), .CO(
        \add_34/carry[8] ), .S(nqp1[7]) );
  HA_X1 \add_34/U1_1_8  ( .A(\add_34/carry[8] ), .B(nq[8]), .CO(
        \add_34/carry[9] ), .S(nqp1[8]) );
  HA_X1 \add_34/U1_1_9  ( .A(\add_34/carry[9] ), .B(nq[9]), .CO(
        \add_34/carry[10] ), .S(nqp1[9]) );
  HA_X1 \add_34/U1_1_10  ( .A(\add_34/carry[10] ), .B(nq[10]), .CO(
        \add_34/carry[11] ), .S(nqp1[10]) );
  HA_X1 \add_34/U1_1_11  ( .A(\add_34/carry[11] ), .B(nq[11]), .CO(
        \add_34/carry[12] ), .S(nqp1[11]) );
  HA_X1 \add_34/U1_1_12  ( .A(\add_34/carry[12] ), .B(nq[12]), .CO(
        \add_34/carry[13] ), .S(nqp1[12]) );
  HA_X1 \add_34/U1_1_13  ( .A(\add_34/carry[13] ), .B(nq[13]), .CO(
        \add_34/carry[14] ), .S(nqp1[13]) );
  HA_X1 \add_34/U1_1_14  ( .A(\add_34/carry[14] ), .B(nq[14]), .CO(
        \add_34/carry[15] ), .S(nqp1[14]) );
  HA_X1 \add_34/U1_1_15  ( .A(\add_34/carry[15] ), .B(nq[15]), .CO(
        \add_34/carry[16] ), .S(nqp1[15]) );
  HA_X1 \add_34/U1_1_16  ( .A(\add_34/carry[16] ), .B(nq[16]), .CO(
        \add_34/carry[17] ), .S(nqp1[16]) );
  HA_X1 \add_34/U1_1_17  ( .A(\add_34/carry[17] ), .B(nq[17]), .CO(
        \add_34/carry[18] ), .S(nqp1[17]) );
  HA_X1 \add_34/U1_1_18  ( .A(\add_34/carry[18] ), .B(nq[18]), .CO(
        \add_34/carry[19] ), .S(nqp1[18]) );
  HA_X1 \add_34/U1_1_19  ( .A(\add_34/carry[19] ), .B(nq[19]), .CO(
        \add_34/carry[20] ), .S(nqp1[19]) );
  HA_X1 \add_34/U1_1_20  ( .A(\add_34/carry[20] ), .B(nq[20]), .CO(
        \add_34/carry[21] ), .S(nqp1[20]) );
  HA_X1 \add_34/U1_1_21  ( .A(\add_34/carry[21] ), .B(nq[21]), .CO(
        \add_34/carry[22] ), .S(nqp1[21]) );
  HA_X1 \add_34/U1_1_22  ( .A(\add_34/carry[22] ), .B(nq[22]), .CO(
        \add_34/carry[23] ), .S(nqp1[22]) );
  HA_X1 \add_34/U1_1_23  ( .A(\add_34/carry[23] ), .B(nq[23]), .CO(
        \add_34/carry[24] ), .S(nqp1[23]) );
  HA_X1 \add_34/U1_1_24  ( .A(\add_34/n2 ), .B(nq[24]), .CO(\add_34/carry[25] ), .S(nqp1[24]) );
  HA_X1 \add_34/U1_1_25  ( .A(\add_34/carry[25] ), .B(nq[25]), .CO(), .S(
        nqp1[25]) );
  HA_X1 \add_34/U1_1_26  ( .A(\add_34/carry[26] ), .B(nq[26]), .CO(
        \add_34/carry[27] ), .S(nqp1[26]) );
  HA_X1 \add_34/U1_1_27  ( .A(\add_34/carry[27] ), .B(nq[27]), .CO(
        \add_34/carry[28] ), .S(nqp1[27]) );
  HA_X1 \add_34/U1_1_29  ( .A(\add_34/carry[29] ), .B(nq[29]), .CO(
        \add_34/carry[30] ), .S(nqp1[29]) );
endmodule

